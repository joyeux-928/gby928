1 1 0 1 0
1 2 0 1 0
1 3 0 1 0
1 4 0 1 0
1 5 0 1 0
1 6 0 1 0
1 7 0 1 0
1 8 0 2 0
1 11 0 2 0
1 14 0 1 0
1 15 0 1 0
1 16 0 2 0
1 19 0 1 0
1 20 0 1 0
1 21 0 1 0
1 22 0 1 0
1 23 0 1 0
1 24 0 1 0
1 25 0 1 0
1 26 0 1 0
1 27 0 1 0
1 28 0 1 0
1 29 0 2 0
1 32 0 1 0
1 33 0 1 0
1 34 0 1 0
1 35 0 1 0
1 36 0 1 0
1 37 0 2 0
1 40 0 2 0
1 43 0 1 0
1 44 0 2 0
1 47 0 1 0
1 48 0 1 0
1 49 0 1 0
1 50 0 1 0
1 51 0 1 0
1 52 0 1 0
1 53 0 1 0
1 54 0 1 0
1 55 0 1 0
1 56 0 1 0
1 57 0 2 0
1 60 0 1 0
1 61 0 1 0
1 62 0 1 0
1 63 0 1 0
1 64 0 1 0
1 65 0 1 0
1 66 0 1 0
1 67 0 1 0
1 68 0 1 0
1 69 0 2 0
1 72 0 1 0
1 73 0 1 0
1 74 0 1 0
1 75 0 1 0
1 76 0 1 0
1 77 0 1 0
1 78 0 1 0
1 79 0 1 0
1 80 0 1 0
1 81 0 1 0
1 82 0 2 0
1 85 0 1 0
1 86 0 1 0
1 87 0 1 0
1 88 0 1 0
1 89 0 1 0
1 90 0 1 0
1 91 0 1 0
1 92 0 1 0
1 93 0 1 0
1 94 0 1 0
1 95 0 1 0
1 96 0 2 0
1 99 0 1 0
1 100 0 1 0
1 101 0 1 0
1 102 0 1 0
1 103 0 1 0
1 104 0 1 0
1 105 0 1 0
1 106 0 1 0
1 107 0 1 0
1 108 0 2 0
1 111 0 1 0
1 112 0 1 0
1 113 0 1 0
1 114 0 1 0
1 115 0 1 0
1 116 0 1 0
1 117 0 1 0
1 118 0 1 0
1 119 0 1 0
1 120 0 2 0
1 123 0 1 0
1 124 0 1 0
1 125 0 1 0
1 126 0 1 0
1 127 0 1 0
1 128 0 1 0
1 129 0 1 0
1 130 0 1 0
1 131 0 1 0
1 132 0 2 0
1 135 0 1 0
1 136 0 1 0
1 137 0 1 0
1 138 0 1 0
1 139 0 1 0
1 140 0 1 0
1 141 0 1 0
1 142 0 1 0
3 143 0 0 0 
3 144 0 0 0 
3 145 0 0 0 
3 146 0 0 0 
3 147 0 0 0 
3 148 0 0 0 
3 149 0 0 0 
3 150 0 0 0 
3 151 0 0 0 
3 152 0 0 0 
3 153 0 0 0 
3 154 0 0 0 
3 155 0 0 0 
3 156 0 0 0 
3 157 0 0 0 
3 158 0 0 0 
3 159 0 0 0 
3 160 0 0 0 
3 161 0 0 0 
3 162 0 0 0 
3 163 0 0 0 
3 164 0 0 0 
3 165 0 0 0 
3 166 0 0 0 
3 167 0 0 0 
3 168 0 0 0 
3 169 0 0 0 
3 170 0 0 0 
3 171 0 0 0 
3 172 0 0 0 
3 173 0 0 0 
3 174 0 0 0 
3 175 0 0 0 
3 176 0 0 0 
3 177 0 0 0 
3 178 0 0 0 
3 179 0 0 0 
3 180 0 0 0 
3 181 0 0 0 
3 182 0 0 0 
3 183 0 0 0 
3 184 0 0 0 
3 185 0 0 0 
3 186 0 0 0 
3 187 0 0 0 
3 188 0 0 0 
3 189 0 0 0 
3 190 0 0 0 
3 191 0 0 0 
3 192 0 0 0 
3 193 0 0 0 
3 194 0 0 0 
3 195 0 0 0 
3 196 0 0 0 
3 197 0 0 0 
3 198 0 0 0 
3 199 0 0 0 
3 200 0 0 0 
3 201 0 0 0 
3 202 0 0 0 
3 203 0 0 0 
3 204 0 0 0 
3 205 0 0 0 
3 206 0 0 0 
3 207 0 0 0 
3 208 0 0 0 
3 209 0 0 0 
3 210 0 0 0 
3 211 0 0 0 
3 212 0 0 0 
3 213 0 0 0 
3 214 0 0 0 
3 215 0 0 0 
3 216 0 0 0 
3 217 0 0 0 
3 218 0 0 0 
1 219 0 4 0
1 224 0 2 0
1 227 0 2 0
1 230 0 1 0
1 231 0 2 0
1 234 0 2 0
1 237 0 3 0
1 241 0 4 0
1 246 0 6 0
1 253 0 2 0
1 256 0 2 0
1 259 0 2 0
1 262 0 1 0
1 263 0 2 0
1 266 0 2 0
1 269 0 2 0
1 272 0 2 0
1 275 0 2 0
1 278 0 2 0
1 281 0 2 0
1 284 0 2 0
1 287 0 2 0
1 290 0 3 0
1 294 0 2 0
1 297 0 3 0
1 301 0 3 0
1 305 0 3 0
1 309 0 3 0
1 313 0 2 0
1 316 0 2 0
1 319 0 2 0
1 322 0 2 0
1 325 0 2 0
1 328 0 2 0
1 331 0 2 0
1 334 0 2 0
1 337 0 2 0
1 340 0 2 0
1 343 0 2 0
1 346 0 2 0
1 349 0 2 0
1 352 0 2 0
1 355 0 2 0
3 398 9 0 1 220
3 400 9 0 1 221
3 401 9 0 1 222
0 405 7 1 2 1 3
0 408 5 1 1 230
3 419 9 0 1 254
3 420 9 0 1 255
0 425 5 1 1 262
3 456 9 0 1 291
3 457 9 0 1 292
3 458 9 0 1 293
0 485 7 1 4 310 306 302 298
0 486 5 1 1 405
3 487 5 0 1 45
3 488 5 0 1 133
3 489 5 0 1 83
3 490 5 0 1 97
3 491 5 0 1 70
3 492 5 0 1 121
3 493 5 0 1 58
3 494 5 0 1 109
0 495 7 1 3 2 15 238
0 496 9 2 1 239
0 499 7 1 2 38 38
0 500 9 2 1 223
0 503 9 2 1 9
0 506 9 2 1 10
0 509 9 11 1 228
0 521 9 11 1 235
0 533 5 3 1 242
0 537 5 5 1 247
0 543 7 1 2 12 248
0 544 7 2 4 134 84 98 46
0 547 7 2 4 122 59 110 71
0 550 9 11 1 229
0 562 9 11 1 236
0 574 5 3 1 257
0 578 5 3 1 260
0 582 9 11 1 320
0 594 9 11 1 323
0 606 5 1 1 329
0 607 5 1 1 332
0 608 5 1 1 335
0 609 5 1 1 338
0 610 5 1 1 341
0 611 5 1 1 344
0 612 5 1 1 353
0 613 9 11 1 321
0 625 9 11 1 324
0 637 9 5 1 17
0 643 9 6 1 18
0 650 5 1 1 356
0 651 7 3 2 7 240
0 655 5 3 1 264
0 659 5 3 1 267
0 663 5 3 1 270
0 667 5 3 1 273
0 671 5 3 1 276
0 675 5 3 1 279
0 679 5 3 1 282
0 683 5 3 1 285
0 687 5 5 1 288
0 693 9 5 1 30
0 699 9 5 1 31
0 705 5 5 1 295
0 711 5 3 1 299
0 715 5 3 1 303
0 719 5 3 1 307
0 723 5 3 1 311
0 727 5 2 1 314
0 730 5 2 1 317
0 733 5 1 1 347
0 734 5 1 1 350
0 735 9 2 1 261
0 738 9 2 1 258
0 741 9 2 1 265
0 744 9 2 1 271
0 747 9 2 1 268
0 750 9 2 1 277
0 753 9 2 1 274
0 756 9 2 1 283
0 759 9 2 1 280
0 762 9 2 1 289
0 765 9 2 1 286
0 768 9 2 1 296
0 771 9 2 1 304
0 774 9 2 1 300
0 777 9 2 1 312
0 780 9 2 1 308
0 783 9 2 1 318
0 786 9 2 1 315
3 792 5 0 1 485
3 799 5 0 1 495
0 800 5 2 1 499
3 805 9 0 1 501
0 900 6 1 2 333 606
0 901 6 1 2 330 607
0 902 6 1 2 339 608
0 903 6 1 2 336 609
0 904 6 1 2 345 610
0 905 6 1 2 342 611
0 998 6 1 2 351 733
0 999 6 1 2 348 734
3 1026 7 0 2 94 502
0 1027 7 1 2 326 652
3 1028 5 0 1 653
3 1029 6 0 2 232 654
0 1032 5 1 1 545
0 1033 5 1 1 548
0 1034 7 2 2 549 546
0 1037 9 4 1 504
0 1042 5 10 1 510
0 1053 5 10 1 522
0 1064 7 1 3 80 511 523
0 1065 7 1 3 68 512 524
0 1066 7 1 3 79 513 525
0 1067 7 1 3 78 514 526
0 1068 7 1 3 77 515 527
0 1069 7 1 2 13 538
0 1070 9 4 1 505
0 1075 5 10 1 551
0 1086 5 10 1 563
0 1097 7 1 3 76 552 564
0 1098 7 1 3 75 553 565
0 1099 7 1 3 74 554 566
0 1100 7 1 3 73 555 567
0 1101 7 1 3 72 556 568
0 1102 5 10 1 583
0 1113 5 10 1 595
0 1124 7 1 3 114 584 596
0 1125 7 1 3 113 585 597
0 1126 7 1 3 112 586 598
0 1127 7 1 3 111 587 599
0 1128 7 1 2 588 600
0 1129 6 3 2 900 901
0 1133 6 3 2 902 903
0 1137 6 2 2 904 905
0 1140 5 1 1 742
0 1141 6 1 2 743 612
0 1142 5 1 1 745
0 1143 5 1 1 748
0 1144 5 1 1 751
0 1145 5 1 1 754
0 1146 5 10 1 614
0 1157 5 10 1 626
0 1168 7 1 3 118 615 627
0 1169 7 1 3 107 616 628
0 1170 7 1 3 117 617 629
0 1171 7 1 3 116 618 630
0 1172 7 1 3 115 619 631
0 1173 5 4 1 638
0 1178 5 5 1 644
0 1184 5 1 1 769
0 1185 6 1 2 770 650
0 1186 5 1 1 772
0 1187 5 1 1 775
0 1188 5 1 1 778
0 1189 5 1 1 781
0 1190 9 4 1 507
0 1195 9 4 1 508
0 1200 5 4 1 694
0 1205 5 4 1 700
0 1210 5 1 1 736
0 1211 5 1 1 739
0 1212 5 1 1 757
0 1213 5 1 1 760
0 1214 5 1 1 763
0 1215 5 1 1 766
0 1216 6 2 2 998 999
0 1219 9 2 1 575
0 1222 9 2 1 579
0 1225 9 2 1 656
0 1228 9 2 1 660
0 1231 9 2 1 664
0 1234 9 2 1 668
0 1237 9 2 1 672
0 1240 9 2 1 676
0 1243 9 2 1 680
0 1246 9 2 1 684
0 1249 5 1 1 784
0 1250 5 1 1 787
0 1251 9 2 1 688
0 1254 9 2 1 706
0 1257 9 2 1 712
0 1260 9 2 1 716
0 1263 9 2 1 720
0 1266 9 2 1 724
3 1269 5 0 1 1027
0 1275 7 1 2 327 1032
0 1276 7 1 2 233 1033
3 1277 9 0 1 1035
0 1302 3 1 2 1069 543
0 1351 6 1 2 354 1140
0 1352 6 1 2 749 1142
0 1353 6 1 2 746 1143
0 1354 6 1 2 755 1144
0 1355 6 1 2 752 1145
0 1395 6 1 2 357 1184
0 1396 6 1 2 776 1186
0 1397 6 1 2 773 1187
0 1398 6 1 2 782 1188
0 1399 6 1 2 779 1189
0 1422 6 1 2 740 1210
0 1423 6 1 2 737 1211
0 1424 6 1 2 761 1212
0 1425 6 1 2 758 1213
0 1426 6 1 2 767 1214
0 1427 6 1 2 764 1215
0 1440 6 1 2 788 1249
0 1441 6 1 2 785 1250
3 1448 5 0 1 1036
0 1449 5 1 1 1275
0 1450 5 1 1 1276
0 1451 7 1 3 93 1043 1054
0 1452 7 1 3 55 516 1055
0 1453 7 1 3 67 1044 528
0 1454 7 1 3 81 1045 1056
0 1455 7 1 3 43 517 1057
0 1456 7 1 3 56 1046 529
0 1457 7 1 3 92 1047 1058
0 1458 7 1 3 54 518 1059
0 1459 7 1 3 66 1048 530
0 1460 7 1 3 91 1049 1060
0 1461 7 1 3 53 519 1061
0 1462 7 1 3 65 1050 531
0 1463 7 1 3 90 1051 1062
0 1464 7 1 3 52 520 1063
0 1465 7 1 3 64 1052 532
0 1466 7 1 3 89 1076 1087
0 1467 7 1 3 51 557 1088
0 1468 7 1 3 63 1077 569
0 1469 7 1 3 88 1078 1089
0 1470 7 1 3 50 558 1090
0 1471 7 1 3 62 1079 570
0 1472 7 1 3 87 1080 1091
0 1473 7 1 3 49 559 1092
0 1474 7 1 2 1081 571
0 1475 7 1 3 86 1082 1093
0 1476 7 1 3 48 560 1094
0 1477 7 1 3 61 1083 572
0 1478 7 1 3 85 1084 1095
0 1479 7 1 3 47 561 1096
0 1480 7 1 3 60 1085 573
0 1481 7 1 3 138 1103 1114
0 1482 7 1 3 102 589 1115
0 1483 7 1 3 126 1104 601
0 1484 7 1 3 137 1105 1116
0 1485 7 1 3 101 590 1117
0 1486 7 1 3 125 1106 602
0 1487 7 1 3 136 1107 1118
0 1488 7 1 3 100 591 1119
0 1489 7 1 3 124 1108 603
0 1490 7 1 3 135 1109 1120
0 1491 7 1 3 99 592 1121
0 1492 7 1 3 123 1110 604
0 1493 7 1 2 1111 1122
0 1494 7 1 2 593 1123
0 1495 7 1 2 1112 605
0 1496 5 2 1 1130
0 1499 5 2 1 1134
0 1502 6 3 2 1351 1141
0 1506 6 3 2 1352 1353
0 1510 6 2 2 1354 1355
0 1513 9 2 1 1138
0 1516 9 2 1 1139
0 1519 5 1 1 1220
0 1520 5 1 1 1223
0 1521 5 1 1 1226
0 1522 5 1 1 1229
0 1523 5 1 1 1232
0 1524 5 1 1 1235
0 1525 5 1 1 1238
0 1526 5 1 1 1241
0 1527 5 1 1 1244
0 1528 5 1 1 1247
0 1529 7 1 3 142 1147 1158
0 1530 7 1 3 106 620 1159
0 1531 7 1 3 130 1148 632
0 1532 7 1 3 131 1149 1160
0 1533 7 1 3 95 621 1161
0 1534 7 1 3 119 1150 633
0 1535 7 1 3 141 1151 1162
0 1536 7 1 3 105 622 1163
0 1537 7 1 3 129 1152 634
0 1538 7 1 3 140 1153 1164
0 1539 7 1 3 104 623 1165
0 1540 7 1 3 128 1154 635
0 1541 7 1 3 139 1155 1166
0 1542 7 1 3 103 624 1167
0 1543 7 1 3 127 1156 636
0 1544 7 1 2 19 1174
0 1545 7 1 2 4 1175
0 1546 7 1 2 20 1176
0 1547 7 1 2 5 1177
0 1548 7 1 2 21 1179
0 1549 7 1 2 22 1180
0 1550 7 1 2 23 1181
0 1551 7 1 2 6 1182
0 1552 7 1 2 24 1183
0 1553 6 3 2 1395 1185
0 1557 6 3 2 1396 1397
0 1561 6 2 2 1398 1399
0 1564 7 1 2 25 1201
0 1565 7 1 2 32 1202
0 1566 7 1 2 26 1203
0 1567 7 1 2 33 1204
0 1568 7 1 2 27 1206
0 1569 7 1 2 34 1207
0 1570 7 1 2 35 1208
0 1571 7 1 2 28 1209
0 1572 5 1 1 1252
0 1573 5 1 1 1255
0 1574 5 1 1 1258
0 1575 5 1 1 1261
0 1576 5 1 1 1264
0 1577 5 1 1 1267
0 1578 6 2 2 1422 1423
0 1581 5 1 1 1217
0 1582 6 2 2 1426 1427
0 1585 6 2 2 1424 1425
0 1588 6 2 2 1440 1441
0 1591 7 4 2 1449 1450
0 1596 3 3 4 1451 1452 1453 1064
0 1600 3 5 4 1454 1455 1456 1065
0 1606 3 5 4 1457 1458 1459 1066
0 1612 3 2 4 1460 1461 1462 1067
0 1615 3 3 4 1463 1464 1465 1068
0 1619 3 4 4 1466 1467 1468 1097
0 1624 3 3 4 1469 1470 1471 1098
0 1628 3 2 4 1472 1473 1474 1099
0 1631 3 2 4 1475 1476 1477 1100
0 1634 3 2 4 1478 1479 1480 1101
0 1637 3 4 4 1481 1482 1483 1124
0 1642 3 4 4 1484 1485 1486 1125
0 1647 3 3 4 1487 1488 1489 1126
0 1651 3 4 4 1490 1491 1492 1127
0 1656 3 3 4 1493 1494 1495 1128
0 1676 3 4 4 1532 1533 1534 1169
0 1681 3 4 4 1535 1536 1537 1170
0 1686 3 3 4 1538 1539 1540 1171
0 1690 3 2 4 1541 1542 1543 1172
0 1708 3 2 4 1529 1530 1531 1168
3 1726 9 0 1 1592
0 1770 5 2 1 1503
0 1773 5 2 1 1507
0 1776 5 1 1 1514
0 1777 5 1 1 1517
0 1778 9 2 1 1511
0 1781 9 2 1 1512
0 1784 7 1 3 1135 1131 1515
0 1785 7 1 3 1500 1497 1518
0 1795 5 2 1 1554
0 1798 5 2 1 1558
0 1801 9 2 1 1562
0 1804 9 2 1 1563
0 1807 5 1 1 1589
0 1808 5 1 1 1579
0 1809 6 1 2 1580 1581
0 1810 5 1 1 1583
0 1811 5 1 1 1586
0 1813 7 1 2 1597 243
0 1814 7 1 2 1607 244
0 1815 7 1 2 1601 245
3 1816 5 0 1 1643
3 1817 5 0 1 1648
3 1818 5 0 1 1638
3 1819 5 0 1 1625
3 1820 5 0 1 1620
3 1821 5 0 1 1616
0 1822 7 1 4 497 225 36 1593
0 1823 7 1 4 498 226 1594 486
0 1824 9 2 1 1598
0 1827 5 2 1 1608
0 1830 7 1 2 1602 539
0 1831 7 1 2 1609 540
0 1832 7 1 2 1621 249
0 1833 5 2 1 1599
0 1836 5 4 1 1603
0 1841 5 6 1 1610
0 1848 9 3 1 1613
0 1852 9 3 1 1617
0 1856 9 6 1 1622
0 1863 9 6 1 1626
0 1870 9 4 1 1629
0 1875 9 4 1 1632
0 1880 9 4 1 1635
0 1885 6 2 2 728 1652
0 1888 6 2 2 731 1657
0 1891 9 2 1 1687
0 1894 7 2 2 1639 425
0 1897 5 2 1 1644
0 1908 7 1 3 1498 1136 1776
0 1909 7 1 3 1132 1501 1777
0 1910 7 1 2 1604 639
0 1911 7 1 2 1611 640
0 1912 7 1 2 1614 641
0 1913 7 1 2 1618 642
0 1914 7 1 2 1623 645
0 1915 7 1 2 1627 646
0 1916 7 1 2 1630 647
0 1917 7 1 2 1633 648
0 1918 7 1 2 1636 649
0 1919 5 1 1 1709
0 1928 7 1 2 1677 695
0 1929 7 1 2 1682 696
0 1930 7 1 2 1688 697
0 1931 7 1 2 1691 698
0 1932 7 1 2 1640 701
0 1933 7 1 2 1645 702
0 1934 7 1 2 1649 703
0 1935 7 1 2 1653 704
0 1936 9 2 1 1605
0 1939 6 1 2 1218 1808
0 1940 6 1 2 1587 1810
0 1941 6 1 2 1584 1811
0 1942 9 2 1 1678
0 1945 9 2 1 1689
0 1948 9 2 1 1683
0 1951 9 2 1 1641
0 1954 9 2 1 1692
0 1957 9 2 1 1650
0 1960 9 2 1 1646
0 1963 9 2 1 1658
0 1966 9 2 1 1654
3 1969 3 0 2 534 1815
3 1970 5 0 1 1822
3 1971 5 0 1 1823
3 2010 9 0 1 1849
3 2012 9 0 1 1853
3 2014 9 0 1 1857
3 2016 9 0 1 1864
3 2018 9 0 1 1871
3 2020 9 0 1 1876
3 2022 9 0 1 1881
0 2028 5 1 1 1779
0 2029 5 1 1 1782
0 2030 4 1 2 1908 1784
0 2031 4 1 2 1909 1785
0 2032 7 1 3 1508 1504 1780
0 2033 7 1 3 1774 1771 1783
0 2034 3 1 2 1571 1935
0 2040 5 1 1 1802
0 2041 5 1 1 1805
0 2042 7 1 3 1559 1555 1803
0 2043 7 1 3 1799 1796 1806
0 2046 6 2 2 1939 1809
0 2049 6 2 2 1940 1941
0 2052 3 2 2 1544 1910
0 2055 3 2 2 1545 1911
0 2058 3 2 2 1546 1912
0 2061 3 2 2 1547 1913
0 2064 3 2 2 1548 1914
0 2067 3 2 2 1549 1915
0 2070 3 2 2 1550 1916
0 2073 3 2 2 1551 1917
0 2076 3 2 2 1552 1918
0 2079 3 2 2 1564 1928
0 2095 3 2 2 1565 1929
0 2098 3 2 2 1566 1930
0 2101 3 2 2 1567 1931
0 2104 3 2 2 1568 1932
0 2107 3 2 2 1569 1933
0 2110 3 2 2 1570 1934
0 2113 7 5 3 1898 1895 41
0 2119 5 1 1 1896
0 2120 6 4 2 408 1828
0 2125 7 1 2 1825 541
0 2126 7 1 2 1854 250
0 2127 7 1 2 1850 542
0 2128 5 6 1 1851
0 2135 5 5 1 1855
0 2141 5 2 1 1865
0 2144 5 2 1 1872
0 2147 5 2 1 1877
0 2150 5 2 1 1882
0 2153 7 1 2 729 1886
0 2154 7 1 2 1887 1655
0 2155 7 1 2 732 1889
0 2156 7 1 2 1890 1659
0 2157 7 1 3 1772 1509 2028
0 2158 7 1 3 1505 1775 2029
0 2171 5 1 1 1943
0 2172 6 1 2 1944 1919
0 2173 5 1 1 1946
0 2174 5 1 1 1949
0 2175 5 1 1 1952
0 2176 5 1 1 1955
0 2177 7 1 3 1797 1560 2040
0 2178 7 1 3 1556 1800 2041
0 2185 9 2 1 1837
0 2188 9 2 1 1834
0 2191 9 2 1 1842
0 2194 5 2 1 1858
0 2197 5 2 1 1829
0 2200 5 1 1 1937
0 2201 9 2 1 1838
0 2204 9 2 1 1835
0 2207 9 2 1 1843
0 2210 9 2 1 1826
0 2213 9 2 1 1844
0 2216 9 2 1 1845
0 2219 6 2 2 2031 2030
0 2234 5 1 1 1958
0 2235 5 1 1 1961
0 2236 5 1 1 1964
0 2237 5 1 1 1967
0 2250 7 2 3 42 1899 2119
0 2266 3 2 2 1831 2126
0 2269 3 2 2 2127 1832
0 2291 3 2 2 2153 2154
0 2294 3 2 2 2155 2156
0 2297 4 1 2 2157 2032
0 2298 4 1 2 2158 2033
0 2300 5 1 1 2047
0 2301 5 1 1 2050
0 2302 6 1 2 2053 1519
0 2303 5 1 1 2054
0 2304 6 1 2 2056 1520
0 2305 5 1 1 2057
0 2306 6 1 2 2059 1521
0 2307 5 1 1 2060
0 2308 6 1 2 2062 1522
0 2309 5 1 1 2063
0 2310 6 1 2 2065 1523
0 2311 5 1 1 2066
0 2312 6 1 2 2068 1524
0 2313 5 1 1 2069
0 2314 6 1 2 2071 1525
0 2315 5 1 1 2072
0 2316 6 1 2 2074 1526
0 2317 5 1 1 2075
0 2318 6 1 2 2077 1527
0 2319 5 1 1 2078
0 2320 6 1 2 2080 1528
0 2321 5 1 1 2081
0 2322 6 1 2 1710 2171
0 2323 6 1 2 1950 2173
0 2324 6 1 2 1947 2174
0 2325 6 1 2 1956 2175
0 2326 6 1 2 1953 2176
0 2327 4 1 2 2177 2042
0 2328 4 1 2 2178 2043
0 2329 6 1 2 2096 1572
0 2330 5 1 1 2097
0 2331 6 1 2 2099 1573
0 2332 5 1 1 2100
0 2333 6 1 2 2102 1574
0 2334 5 1 1 2103
0 2335 6 1 2 2105 1575
0 2336 5 1 1 2106
0 2337 6 1 2 2108 1576
0 2338 5 1 1 2109
0 2339 6 1 2 2111 1577
0 2340 5 1 1 2112
0 2354 6 1 2 1962 2234
0 2355 6 1 2 1959 2235
0 2356 6 1 2 1968 2236
0 2357 6 1 2 1965 2237
0 2358 7 1 2 2121 535
0 2359 5 2 1 2114
0 2364 5 1 1 2186
0 2365 5 1 1 2189
0 2366 5 1 1 2192
0 2367 5 1 1 2195
0 2368 9 3 1 2122
0 2372 5 1 1 2202
0 2373 5 1 1 2205
0 2374 5 1 1 2208
0 2375 5 1 1 2211
0 2376 5 1 1 2214
0 2377 5 4 1 2115
0 2382 9 3 1 2116
0 2386 7 1 2 2123 251
3 2387 9 0 1 2267
3 2388 9 0 1 2268
3 2389 9 0 1 2270
3 2390 9 0 1 2271
0 2391 9 3 1 2117
0 2395 5 4 1 2118
0 2400 6 1 2 2220 2300
0 2403 5 1 1 2217
0 2406 5 1 1 2221
0 2407 6 1 2 1221 2303
0 2408 6 1 2 1224 2305
0 2409 6 1 2 1227 2307
0 2410 6 1 2 1230 2309
0 2411 6 1 2 1233 2311
0 2412 6 1 2 1236 2313
0 2413 6 1 2 1239 2315
0 2414 6 1 2 1242 2317
0 2415 6 1 2 1245 2319
0 2416 6 1 2 1248 2321
0 2417 6 3 2 2322 2172
0 2421 6 3 2 2323 2324
0 2425 6 2 2 2325 2326
0 2428 6 1 2 1253 2330
0 2429 6 1 2 1256 2332
0 2430 6 1 2 1259 2334
0 2431 6 1 2 1262 2336
0 2432 6 1 2 1265 2338
0 2433 6 1 2 1268 2340
0 2434 9 2 1 2129
0 2437 9 2 1 2136
0 2440 9 2 1 2145
0 2443 9 2 1 2142
0 2446 9 2 1 2151
0 2449 9 2 1 2148
0 2452 5 1 1 2198
0 2453 6 1 2 2199 2200
0 2454 9 2 1 2130
0 2457 9 2 1 2146
0 2460 9 2 1 2143
0 2463 9 2 1 2152
0 2466 9 2 1 2149
0 2469 5 2 1 2124
0 2472 9 2 1 2131
0 2475 9 2 1 2137
0 2478 9 2 1 2132
0 2481 9 2 1 2138
0 2484 6 2 2 2298 2297
0 2487 6 2 2 2356 2357
0 2490 6 2 2 2354 2355
0 2493 6 2 2 2328 2327
3 2496 3 0 2 2358 1814
0 2503 6 1 2 2190 2364
0 2504 6 1 2 2187 2365
0 2510 6 1 2 2206 2372
0 2511 6 1 2 2203 2373
0 2521 3 2 2 1830 2386
0 2528 6 1 2 2048 2406
0 2531 5 2 1 2292
0 2534 5 2 1 2295
0 2537 9 2 1 2251
0 2540 9 2 1 2252
0 2544 6 1 2 2302 2407
0 2545 6 1 2 2304 2408
0 2546 6 1 2 2306 2409
0 2547 6 1 2 2308 2410
0 2548 6 1 2 2310 2411
0 2549 6 1 2 2312 2412
0 2550 6 1 2 2314 2413
0 2551 6 1 2 2316 2414
0 2552 6 1 2 2318 2415
0 2553 6 1 2 2320 2416
0 2563 6 1 2 2329 2428
0 2564 6 1 2 2331 2429
0 2565 6 1 2 2333 2430
0 2566 6 1 2 2335 2431
0 2567 6 1 2 2337 2432
0 2568 6 1 2 2339 2433
0 2579 6 1 2 1938 2452
0 2603 9 3 1 2360
0 2607 7 1 2 1883 2378
0 2608 7 1 2 1679 2379
0 2609 7 1 2 1684 2380
0 2610 7 1 2 1892 2381
0 2611 7 1 2 1859 2383
0 2612 7 1 2 1866 2384
0 2613 6 3 2 2503 2504
0 2617 5 1 1 2435
0 2618 6 1 2 2436 2366
0 2619 6 1 2 2438 2367
0 2620 5 1 1 2439
0 2621 5 2 1 2369
0 2624 6 3 2 2510 2511
0 2628 5 1 1 2455
0 2629 6 1 2 2456 2374
0 2630 5 1 1 2473
0 2631 7 1 2 1860 2392
0 2632 7 1 2 1867 2393
0 2633 7 1 2 1884 2396
0 2634 7 1 2 1680 2397
0 2635 7 1 2 1685 2398
0 2636 7 1 2 1893 2399
0 2638 5 4 1 2385
3 2643 9 0 1 2522
3 2644 9 0 1 2523
0 2645 5 1 1 2476
0 2646 5 4 1 2394
0 2652 6 1 2 2528 2400
0 2655 5 1 1 2479
0 2656 5 1 1 2482
0 2659 9 3 1 2361
0 2663 5 1 1 2485
0 2664 6 1 2 2486 2301
0 2665 5 1 1 2553
0 2666 5 1 1 2552
0 2667 5 1 1 2551
0 2668 5 1 1 2550
0 2669 5 1 1 2549
0 2670 5 1 1 2548
0 2671 5 1 1 2547
0 2672 5 1 1 2546
0 2673 5 1 1 2545
0 2674 5 1 1 2544
0 2675 5 1 1 2568
0 2676 5 1 1 2567
0 2677 5 1 1 2566
0 2678 5 1 1 2565
0 2679 5 1 1 2564
0 2680 5 1 1 2563
0 2681 5 2 1 2418
0 2684 5 2 1 2422
0 2687 9 2 1 2426
0 2690 9 2 1 2427
0 2693 5 1 1 2494
0 2694 6 1 2 2495 1807
0 2695 5 1 1 2441
0 2696 5 1 1 2444
0 2697 5 1 1 2447
0 2698 5 1 1 2450
0 2699 5 1 1 2458
0 2700 5 1 1 2461
0 2701 5 1 1 2464
0 2702 5 1 1 2467
0 2703 6 2 2 2579 2453
0 2706 5 1 1 2470
0 2707 5 1 1 2488
0 2708 5 1 1 2491
0 2709 7 1 2 2296 2535
0 2710 7 1 2 2293 2532
0 2719 6 1 2 2193 2617
0 2720 6 1 2 2196 2620
0 2726 6 1 2 2209 2628
0 2729 9 4 1 2538
0 2738 9 4 1 2539
0 2743 5 1 1 2652
0 2747 6 1 2 2051 2663
0 2748 7 1 5 2665 2666 2667 2668 2669
0 2749 7 1 5 2670 2671 2672 2673 2674
0 2750 7 1 2 2034 2675
0 2751 7 1 5 2676 2677 2678 2679 2680
0 2760 6 1 2 1590 2693
0 2761 9 4 1 2541
0 2766 9 4 1 2542
0 2771 6 1 2 2445 2695
0 2772 6 1 2 2442 2696
0 2773 6 1 2 2451 2697
0 2774 6 1 2 2448 2698
0 2775 6 1 2 2462 2699
0 2776 6 1 2 2459 2700
0 2777 6 1 2 2468 2701
0 2778 6 1 2 2465 2702
0 2781 6 1 2 2492 2707
0 2782 6 1 2 2489 2708
0 2783 3 1 2 2709 2536
0 2784 3 1 2 2710 2533
0 2789 7 1 2 1861 2639
0 2790 7 1 2 1868 2640
0 2791 7 1 2 1873 2641
0 2792 7 1 2 1878 2642
0 2793 5 2 1 2614
0 2796 6 3 2 2719 2618
0 2800 6 2 2 2619 2720
0 2803 5 2 1 2625
0 2806 6 2 2 2726 2629
0 2809 7 1 2 1862 2647
0 2810 7 1 2 1869 2648
0 2811 7 1 2 1874 2649
0 2812 7 1 2 1879 2650
0 2817 7 2 2 2743 14
0 2820 9 5 1 2604
0 2826 6 2 2 2747 2664
0 2829 7 1 2 2748 2749
0 2830 7 1 2 2750 2751
0 2831 9 5 1 2660
0 2837 5 1 1 2688
0 2838 5 1 1 2691
0 2839 7 1 3 2423 2419 2689
0 2840 7 1 3 2685 2682 2692
0 2841 6 2 2 2760 2694
0 2844 9 5 1 2605
0 2854 9 4 1 2606
0 2859 9 5 1 2661
0 2869 9 4 1 2662
0 2874 6 2 2 2773 2774
0 2877 6 2 2 2771 2772
0 2880 5 1 1 2704
0 2881 6 1 2 2705 2706
0 2882 6 2 2 2777 2778
0 2885 6 2 2 2775 2776
0 2888 6 2 2 2781 2782
3 2891 6 0 2 2783 2784
0 2894 7 1 2 2607 2730
0 2895 7 1 2 2608 2731
0 2896 7 1 2 2609 2732
0 2897 7 1 2 2610 2733
0 2898 3 1 2 2789 2611
0 2899 3 1 2 2790 2612
0 2900 7 1 2 2791 1038
0 2901 7 1 2 2792 1039
0 2914 3 1 2 2809 2631
0 2915 3 1 2 2810 2632
0 2916 7 1 2 2811 1071
0 2917 7 1 2 2812 1072
0 2918 7 1 2 2633 2739
0 2919 7 1 2 2634 2740
0 2920 7 1 2 2635 2741
0 2921 7 1 2 2636 2742
3 2925 9 0 1 2818
0 2931 7 2 3 2829 2830 1302
0 2938 7 1 3 2683 2424 2837
0 2939 7 1 3 2420 2686 2838
0 2963 6 1 2 2471 2880
3 2970 5 0 1 2842
3 2971 5 0 1 2827
0 2972 5 2 1 2894
0 2975 5 2 1 2895
0 2978 5 2 1 2896
0 2981 5 2 1 2897
0 2984 7 1 2 2898 1040
0 2985 7 1 2 2899 1041
0 2986 5 2 1 2900
0 2989 5 2 1 2901
0 2992 5 2 1 2797
0 2995 9 2 1 2801
0 2998 9 2 1 2802
0 3001 9 2 1 2807
0 3004 9 2 1 2808
0 3007 7 1 2 576 2821
0 3008 7 1 2 2914 1073
0 3009 7 1 2 2915 1074
0 3010 5 2 1 2916
0 3013 5 2 1 2917
0 3016 5 2 1 2918
0 3019 5 2 1 2919
0 3022 5 2 1 2920
0 3025 5 2 1 2921
0 3028 5 1 1 2819
0 3029 7 1 2 577 2832
0 3030 5 4 1 2822
0 3035 7 1 2 580 2823
0 3036 7 1 2 657 2824
0 3037 7 1 2 661 2825
3 3038 9 0 1 2932
0 3039 5 4 1 2833
0 3044 7 1 2 581 2834
0 3045 7 1 2 658 2835
0 3046 7 1 2 662 2836
0 3047 4 1 2 2938 2839
0 3048 4 1 2 2939 2840
0 3049 5 1 1 2889
0 3050 5 2 1 2845
0 3053 7 1 2 665 2846
0 3054 7 1 2 669 2847
0 3055 7 1 2 673 2848
0 3056 7 1 2 677 2849
0 3057 7 1 2 681 2855
0 3058 7 1 2 685 2856
0 3059 7 1 2 689 2857
0 3060 7 1 2 707 2858
0 3061 5 2 1 2860
0 3064 7 1 2 666 2861
0 3065 7 1 2 670 2862
0 3066 7 1 2 674 2863
0 3067 7 1 2 678 2864
0 3068 7 1 2 682 2870
0 3069 7 1 2 686 2871
0 3070 7 1 2 690 2872
0 3071 7 1 2 708 2873
0 3072 5 1 1 2875
0 3073 5 1 1 2878
0 3074 5 1 1 2883
0 3075 5 1 1 2886
0 3076 6 2 2 2881 2963
3 3079 5 0 1 2933
0 3088 5 2 1 2984
0 3091 5 2 1 2985
0 3110 5 2 1 3008
0 3113 5 2 1 3009
0 3137 7 2 2 3055 1191
0 3140 7 2 2 3056 1192
0 3143 7 2 2 3057 2762
0 3146 7 2 2 3058 2763
0 3149 7 2 2 3059 2764
0 3152 7 2 2 3060 2765
0 3157 7 2 2 3066 1196
0 3160 7 2 2 3067 1197
0 3163 7 2 2 3068 2767
0 3166 7 2 2 3069 2768
0 3169 7 2 2 3070 2769
0 3172 7 2 2 3071 2770
0 3175 6 1 2 2879 3072
0 3176 6 1 2 2876 3073
0 3177 6 1 2 2887 3074
0 3178 6 1 2 2884 3075
0 3180 6 2 2 3048 3047
0 3187 5 1 1 2996
0 3188 5 1 1 2999
0 3189 5 1 1 3002
0 3190 5 1 1 3005
0 3191 7 1 3 2798 2615 2997
0 3192 7 1 3 2993 2794 3000
0 3193 7 1 3 2626 2370 3003
0 3194 7 1 3 2804 2622 3006
0 3195 6 1 2 3077 2375
0 3196 5 1 1 3078
0 3197 7 1 2 691 3031
0 3208 7 1 2 692 3040
0 3215 7 1 2 709 3032
0 3216 7 1 2 713 3033
0 3217 7 1 2 717 3034
0 3218 7 1 2 710 3041
0 3219 7 1 2 714 3042
0 3220 7 1 2 718 3043
0 3222 7 1 2 721 3051
0 3223 7 1 2 725 3052
0 3230 7 1 2 722 3062
0 3231 7 1 2 726 3063
0 3238 6 2 2 3175 3176
0 3241 6 2 2 3177 3178
0 3244 9 2 1 2982
0 3247 9 2 1 2979
0 3250 9 2 1 2976
0 3253 9 2 1 2973
0 3256 9 2 1 2990
0 3259 9 2 1 2987
0 3262 9 2 1 3026
0 3265 9 2 1 3023
0 3268 9 2 1 3020
0 3271 9 2 1 3017
0 3274 9 2 1 3014
0 3277 9 2 1 3011
0 3281 7 1 3 2795 2799 3187
0 3282 7 1 3 2616 2994 3188
0 3283 7 1 3 2623 2627 3189
0 3284 7 1 3 2371 2805 3190
0 3286 6 1 2 2212 3196
0 3288 3 1 2 3197 3007
0 3289 6 1 2 3181 3049
0 3291 7 1 2 3153 2983
0 3293 7 1 2 3150 2980
0 3295 7 1 2 3147 2977
0 3296 7 1 2 2974 3144
0 3299 7 1 2 3141 2991
0 3301 7 1 2 3138 2988
0 3302 3 1 2 3208 3029
0 3304 7 1 2 3173 3027
0 3306 7 1 2 3170 3024
0 3308 7 1 2 3167 3021
0 3309 7 1 2 3018 3164
0 3312 7 1 2 3161 3015
0 3314 7 1 2 3158 3012
0 3315 3 2 2 3215 3035
0 3318 3 2 2 3216 3036
0 3321 3 2 2 3217 3037
0 3324 3 2 2 3218 3044
0 3327 3 2 2 3219 3045
0 3330 3 2 2 3220 3046
0 3333 5 1 1 3182
0 3334 3 1 2 3222 3053
0 3335 3 1 2 3223 3054
0 3336 3 1 2 3230 3064
0 3337 3 1 2 3231 3065
0 3340 9 2 1 3154
0 3344 9 2 1 3151
0 3348 9 2 1 3148
0 3352 9 2 1 3145
0 3356 9 2 1 3142
0 3360 9 2 1 3139
0 3364 9 2 1 3092
0 3367 9 2 1 3089
0 3370 9 2 1 3174
0 3374 9 2 1 3171
0 3378 9 2 1 3168
0 3382 9 2 1 3165
0 3386 9 2 1 3162
0 3390 9 2 1 3159
0 3394 9 2 1 3114
0 3397 9 2 1 3111
0 3400 6 1 2 3195 3286
0 3401 4 1 2 3281 3191
0 3402 4 1 2 3282 3192
0 3403 4 1 2 3283 3193
0 3404 4 1 2 3284 3194
0 3405 5 1 1 3239
0 3406 5 1 1 3242
0 3409 7 1 2 3288 1839
0 3410 6 1 2 2890 3333
0 3412 5 1 1 3245
0 3414 5 1 1 3248
0 3416 5 1 1 3251
0 3418 5 1 1 3254
0 3420 5 1 1 3257
0 3422 5 1 1 3260
0 3428 7 1 2 3302 1840
0 3430 5 1 1 3263
0 3432 5 1 1 3266
0 3434 5 1 1 3269
0 3436 5 1 1 3272
0 3438 5 1 1 3275
0 3440 5 1 1 3278
0 3450 7 2 2 3334 1193
0 3453 7 2 2 3335 1194
0 3456 7 2 2 3336 1198
0 3459 7 2 2 3337 1199
0 3478 7 1 2 3400 536
0 3479 7 1 2 3319 2133
0 3480 7 1 2 3316 1846
0 3481 6 1 2 3410 3289
0 3482 5 1 1 3341
0 3483 6 1 2 3342 3412
0 3484 5 1 1 3345
0 3485 6 1 2 3346 3414
0 3486 5 1 1 3349
0 3487 6 1 2 3350 3416
0 3488 5 1 1 3353
0 3489 6 1 2 3354 3418
0 3490 5 1 1 3357
0 3491 6 1 2 3358 3420
0 3492 5 1 1 3361
0 3493 6 1 2 3362 3422
0 3494 5 1 1 3365
0 3496 5 1 1 3368
0 3498 7 1 2 3322 2139
0 3499 7 1 2 3328 2134
0 3500 7 1 2 3325 1847
0 3501 5 1 1 3371
0 3502 6 1 2 3372 3430
0 3503 5 1 1 3375
0 3504 6 1 2 3376 3432
0 3505 5 1 1 3379
0 3506 6 1 2 3380 3434
0 3507 5 1 1 3383
0 3508 6 1 2 3384 3436
0 3509 5 1 1 3387
0 3510 6 1 2 3388 3438
0 3511 5 1 1 3391
0 3512 6 1 2 3392 3440
0 3513 5 1 1 3395
0 3515 5 1 1 3398
0 3517 7 1 2 3331 2140
0 3522 6 2 2 3402 3401
0 3525 6 2 2 3404 3403
0 3528 9 2 1 3320
0 3531 9 2 1 3317
0 3534 9 2 1 3323
0 3537 9 2 1 3329
0 3540 9 2 1 3326
0 3543 9 2 1 3332
3 3546 3 0 2 3478 1813
0 3551 5 1 1 3481
0 3552 6 1 2 3246 3482
0 3553 6 1 2 3249 3484
0 3554 6 1 2 3252 3486
0 3555 6 1 2 3255 3488
0 3556 6 1 2 3258 3490
0 3557 6 1 2 3261 3492
0 3558 7 1 2 3454 3093
0 3559 7 1 2 3451 3090
0 3563 6 1 2 3264 3501
0 3564 6 1 2 3267 3503
0 3565 6 1 2 3270 3505
0 3566 6 1 2 3273 3507
0 3567 6 1 2 3276 3509
0 3568 6 1 2 3279 3511
0 3569 7 1 2 3460 3115
0 3570 7 1 2 3457 3112
0 3576 9 2 1 3455
0 3579 9 2 1 3452
0 3585 9 2 1 3461
0 3588 9 2 1 3458
0 3592 5 1 1 3523
0 3593 6 1 2 3524 3405
0 3594 5 1 1 3526
0 3595 6 1 2 3527 3406
0 3596 5 1 1 3529
0 3597 6 1 2 3530 2630
0 3598 6 1 2 3532 2376
0 3599 5 1 1 3533
0 3600 7 2 2 3551 801
0 3603 6 4 2 3552 3483
0 3608 6 3 2 3553 3485
0 3612 6 2 2 3554 3487
0 3615 6 1 2 3555 3489
0 3616 6 5 2 3556 3491
0 3622 6 4 2 3557 3493
0 3629 5 1 1 3535
0 3630 6 1 2 3536 2645
0 3631 5 1 1 3538
0 3632 6 1 2 3539 2655
0 3633 6 1 2 3541 2403
0 3634 5 1 1 3542
0 3635 6 4 2 3563 3502
0 3640 6 3 2 3564 3504
0 3644 6 2 2 3565 3506
0 3647 6 1 2 3566 3508
0 3648 6 5 2 3567 3510
0 3654 6 4 2 3568 3512
0 3661 5 1 1 3544
0 3662 6 1 2 3545 2656
0 3667 6 1 2 3240 3592
0 3668 6 1 2 3243 3594
0 3669 6 1 2 2474 3596
0 3670 6 1 2 2215 3599
3 3671 9 0 1 3601
0 3691 5 1 1 3577
0 3692 6 1 2 3578 3494
0 3693 5 1 1 3580
0 3694 6 1 2 3581 3496
0 3695 6 1 2 2477 3629
0 3696 6 1 2 2480 3631
0 3697 6 1 2 2218 3634
0 3716 5 1 1 3586
0 3717 6 1 2 3587 3513
0 3718 5 1 1 3589
0 3719 6 1 2 3590 3515
0 3720 6 1 2 2483 3661
0 3721 6 1 2 3667 3593
0 3722 6 1 2 3668 3595
0 3723 6 2 2 3669 3597
0 3726 6 1 2 3670 3598
0 3727 5 1 1 3602
0 3728 6 1 2 3366 3691
0 3729 6 1 2 3369 3693
0 3730 6 1 2 3695 3630
0 3731 7 1 4 3609 3615 3613 3604
0 3732 7 1 2 3605 3293
0 3733 7 1 3 3610 3606 3295
0 3734 7 1 4 3614 3607 3296 3611
0 3735 7 1 2 3617 3301
0 3736 7 1 3 3623 3618 3558
0 3737 6 2 2 3696 3632
0 3740 6 1 2 3697 3633
0 3741 6 1 2 3396 3716
0 3742 6 1 2 3399 3718
0 3743 6 1 2 3720 3662
0 3744 7 1 4 3641 3647 3645 3636
0 3745 7 1 2 3637 3306
0 3746 7 1 3 3642 3638 3308
0 3747 7 1 4 3646 3639 3309 3643
0 3748 7 1 2 3649 3314
0 3749 7 1 3 3655 3650 3569
0 3750 5 1 1 3721
0 3753 7 1 2 3722 252
0 3754 6 3 2 3728 3692
0 3758 6 2 2 3729 3694
0 3761 5 1 1 3731
0 3762 3 2 4 3291 3732 3733 3734
0 3767 6 3 2 3741 3717
0 3771 6 2 2 3742 3719
0 3774 5 1 1 3744
0 3775 3 2 4 3304 3745 3746 3747
0 3778 7 1 2 3724 3480
0 3779 7 1 3 3726 3725 3409
0 3780 3 2 2 2125 3753
0 3790 7 2 2 3750 802
0 3793 7 1 2 3738 3500
0 3794 7 1 3 3740 3739 3428
0 3802 3 1 3 3479 3778 3779
3 3803 9 0 1 3781
3 3804 9 0 1 3782
0 3805 5 1 1 3763
0 3806 7 1 5 3624 3730 3755 3619 3759
0 3807 7 1 4 3756 3620 3559 3625
0 3808 7 1 5 3760 3757 3621 3498 3626
3 3809 9 0 1 3791
0 3811 3 1 3 3499 3793 3794
0 3812 5 1 1 3776
0 3813 7 1 5 3656 3743 3768 3651 3772
0 3814 7 1 4 3769 3652 3570 3657
0 3815 7 1 5 3773 3770 3653 3517 3658
0 3816 3 1 5 3299 3735 3736 3807 3808
0 3817 7 1 2 3806 3802
0 3818 6 1 2 3805 3761
0 3819 5 1 1 3792
0 3820 3 1 5 3312 3748 3749 3814 3815
0 3821 7 1 2 3813 3811
0 3822 6 1 2 3812 3774
0 3823 3 2 2 3816 3817
0 3826 7 1 3 3727 3819 2843
0 3827 3 2 2 3820 3821
0 3834 5 1 1 3824
0 3835 7 1 2 3818 3825
0 3836 5 1 1 3828
0 3837 7 1 2 3822 3829
0 3838 7 1 2 3764 3834
0 3839 7 1 2 3777 3836
0 3840 3 2 2 3838 3835
0 3843 3 3 2 3839 3837
3 3851 9 0 1 3844
0 3852 6 2 2 3845 3841
0 3857 7 1 2 3846 3853
0 3858 7 1 2 3854 3842
0 3859 3 2 2 3857 3858
0 3864 5 2 1 3860
0 3869 7 1 2 3861 3865
0 3870 3 2 2 3869 3866
3 3875 5 0 1 3871
0 3876 7 1 3 2828 3028 3872
0 3877 7 2 3 3826 3876 1595
3 3881 9 0 1 3878
3 3882 5 0 1 3879
2 9 1 8
2 10 1 8
2 12 1 11
2 13 1 11
2 17 1 16
2 18 1 16
2 30 1 29
2 31 1 29
2 38 1 37
2 39 1 37
2 41 1 40
2 42 1 40
2 45 1 44
2 46 1 44
2 58 1 57
2 59 1 57
2 70 1 69
2 71 1 69
2 83 1 82
2 84 1 82
2 97 1 96
2 98 1 96
2 109 1 108
2 110 1 108
2 121 1 120
2 122 1 120
2 133 1 132
2 134 1 132
2 220 1 219
2 221 1 219
2 222 1 219
2 223 1 219
2 225 1 224
2 226 1 224
2 228 1 227
2 229 1 227
2 232 1 231
2 233 1 231
2 235 1 234
2 236 1 234
2 238 1 237
2 239 1 237
2 240 1 237
2 242 1 241
2 243 1 241
2 244 1 241
2 245 1 241
2 247 1 246
2 248 1 246
2 249 1 246
2 250 1 246
2 251 1 246
2 252 1 246
2 254 1 253
2 255 1 253
2 257 1 256
2 258 1 256
2 260 1 259
2 261 1 259
2 264 1 263
2 265 1 263
2 267 1 266
2 268 1 266
2 270 1 269
2 271 1 269
2 273 1 272
2 274 1 272
2 276 1 275
2 277 1 275
2 279 1 278
2 280 1 278
2 282 1 281
2 283 1 281
2 285 1 284
2 286 1 284
2 288 1 287
2 289 1 287
2 291 1 290
2 292 1 290
2 293 1 290
2 295 1 294
2 296 1 294
2 298 1 297
2 299 1 297
2 300 1 297
2 302 1 301
2 303 1 301
2 304 1 301
2 306 1 305
2 307 1 305
2 308 1 305
2 310 1 309
2 311 1 309
2 312 1 309
2 314 1 313
2 315 1 313
2 317 1 316
2 318 1 316
2 320 1 319
2 321 1 319
2 323 1 322
2 324 1 322
2 326 1 325
2 327 1 325
2 329 1 328
2 330 1 328
2 332 1 331
2 333 1 331
2 335 1 334
2 336 1 334
2 338 1 337
2 339 1 337
2 341 1 340
2 342 1 340
2 344 1 343
2 345 1 343
2 347 1 346
2 348 1 346
2 350 1 349
2 351 1 349
2 353 1 352
2 354 1 352
2 356 1 355
2 357 1 355
2 497 1 496
2 498 1 496
2 501 1 500
2 502 1 500
2 504 1 503
2 505 1 503
2 507 1 506
2 508 1 506
2 510 1 509
2 511 1 509
2 512 1 509
2 513 1 509
2 514 1 509
2 515 1 509
2 516 1 509
2 517 1 509
2 518 1 509
2 519 1 509
2 520 1 509
2 522 1 521
2 523 1 521
2 524 1 521
2 525 1 521
2 526 1 521
2 527 1 521
2 528 1 521
2 529 1 521
2 530 1 521
2 531 1 521
2 532 1 521
2 534 1 533
2 535 1 533
2 536 1 533
2 538 1 537
2 539 1 537
2 540 1 537
2 541 1 537
2 542 1 537
2 545 1 544
2 546 1 544
2 548 1 547
2 549 1 547
2 551 1 550
2 552 1 550
2 553 1 550
2 554 1 550
2 555 1 550
2 556 1 550
2 557 1 550
2 558 1 550
2 559 1 550
2 560 1 550
2 561 1 550
2 563 1 562
2 564 1 562
2 565 1 562
2 566 1 562
2 567 1 562
2 568 1 562
2 569 1 562
2 570 1 562
2 571 1 562
2 572 1 562
2 573 1 562
2 575 1 574
2 576 1 574
2 577 1 574
2 579 1 578
2 580 1 578
2 581 1 578
2 583 1 582
2 584 1 582
2 585 1 582
2 586 1 582
2 587 1 582
2 588 1 582
2 589 1 582
2 590 1 582
2 591 1 582
2 592 1 582
2 593 1 582
2 595 1 594
2 596 1 594
2 597 1 594
2 598 1 594
2 599 1 594
2 600 1 594
2 601 1 594
2 602 1 594
2 603 1 594
2 604 1 594
2 605 1 594
2 614 1 613
2 615 1 613
2 616 1 613
2 617 1 613
2 618 1 613
2 619 1 613
2 620 1 613
2 621 1 613
2 622 1 613
2 623 1 613
2 624 1 613
2 626 1 625
2 627 1 625
2 628 1 625
2 629 1 625
2 630 1 625
2 631 1 625
2 632 1 625
2 633 1 625
2 634 1 625
2 635 1 625
2 636 1 625
2 638 1 637
2 639 1 637
2 640 1 637
2 641 1 637
2 642 1 637
2 644 1 643
2 645 1 643
2 646 1 643
2 647 1 643
2 648 1 643
2 649 1 643
2 652 1 651
2 653 1 651
2 654 1 651
2 656 1 655
2 657 1 655
2 658 1 655
2 660 1 659
2 661 1 659
2 662 1 659
2 664 1 663
2 665 1 663
2 666 1 663
2 668 1 667
2 669 1 667
2 670 1 667
2 672 1 671
2 673 1 671
2 674 1 671
2 676 1 675
2 677 1 675
2 678 1 675
2 680 1 679
2 681 1 679
2 682 1 679
2 684 1 683
2 685 1 683
2 686 1 683
2 688 1 687
2 689 1 687
2 690 1 687
2 691 1 687
2 692 1 687
2 694 1 693
2 695 1 693
2 696 1 693
2 697 1 693
2 698 1 693
2 700 1 699
2 701 1 699
2 702 1 699
2 703 1 699
2 704 1 699
2 706 1 705
2 707 1 705
2 708 1 705
2 709 1 705
2 710 1 705
2 712 1 711
2 713 1 711
2 714 1 711
2 716 1 715
2 717 1 715
2 718 1 715
2 720 1 719
2 721 1 719
2 722 1 719
2 724 1 723
2 725 1 723
2 726 1 723
2 728 1 727
2 729 1 727
2 731 1 730
2 732 1 730
2 736 1 735
2 737 1 735
2 739 1 738
2 740 1 738
2 742 1 741
2 743 1 741
2 745 1 744
2 746 1 744
2 748 1 747
2 749 1 747
2 751 1 750
2 752 1 750
2 754 1 753
2 755 1 753
2 757 1 756
2 758 1 756
2 760 1 759
2 761 1 759
2 763 1 762
2 764 1 762
2 766 1 765
2 767 1 765
2 769 1 768
2 770 1 768
2 772 1 771
2 773 1 771
2 775 1 774
2 776 1 774
2 778 1 777
2 779 1 777
2 781 1 780
2 782 1 780
2 784 1 783
2 785 1 783
2 787 1 786
2 788 1 786
2 801 1 800
2 802 1 800
2 1035 1 1034
2 1036 1 1034
2 1038 1 1037
2 1039 1 1037
2 1040 1 1037
2 1041 1 1037
2 1043 1 1042
2 1044 1 1042
2 1045 1 1042
2 1046 1 1042
2 1047 1 1042
2 1048 1 1042
2 1049 1 1042
2 1050 1 1042
2 1051 1 1042
2 1052 1 1042
2 1054 1 1053
2 1055 1 1053
2 1056 1 1053
2 1057 1 1053
2 1058 1 1053
2 1059 1 1053
2 1060 1 1053
2 1061 1 1053
2 1062 1 1053
2 1063 1 1053
2 1071 1 1070
2 1072 1 1070
2 1073 1 1070
2 1074 1 1070
2 1076 1 1075
2 1077 1 1075
2 1078 1 1075
2 1079 1 1075
2 1080 1 1075
2 1081 1 1075
2 1082 1 1075
2 1083 1 1075
2 1084 1 1075
2 1085 1 1075
2 1087 1 1086
2 1088 1 1086
2 1089 1 1086
2 1090 1 1086
2 1091 1 1086
2 1092 1 1086
2 1093 1 1086
2 1094 1 1086
2 1095 1 1086
2 1096 1 1086
2 1103 1 1102
2 1104 1 1102
2 1105 1 1102
2 1106 1 1102
2 1107 1 1102
2 1108 1 1102
2 1109 1 1102
2 1110 1 1102
2 1111 1 1102
2 1112 1 1102
2 1114 1 1113
2 1115 1 1113
2 1116 1 1113
2 1117 1 1113
2 1118 1 1113
2 1119 1 1113
2 1120 1 1113
2 1121 1 1113
2 1122 1 1113
2 1123 1 1113
2 1130 1 1129
2 1131 1 1129
2 1132 1 1129
2 1134 1 1133
2 1135 1 1133
2 1136 1 1133
2 1138 1 1137
2 1139 1 1137
2 1147 1 1146
2 1148 1 1146
2 1149 1 1146
2 1150 1 1146
2 1151 1 1146
2 1152 1 1146
2 1153 1 1146
2 1154 1 1146
2 1155 1 1146
2 1156 1 1146
2 1158 1 1157
2 1159 1 1157
2 1160 1 1157
2 1161 1 1157
2 1162 1 1157
2 1163 1 1157
2 1164 1 1157
2 1165 1 1157
2 1166 1 1157
2 1167 1 1157
2 1174 1 1173
2 1175 1 1173
2 1176 1 1173
2 1177 1 1173
2 1179 1 1178
2 1180 1 1178
2 1181 1 1178
2 1182 1 1178
2 1183 1 1178
2 1191 1 1190
2 1192 1 1190
2 1193 1 1190
2 1194 1 1190
2 1196 1 1195
2 1197 1 1195
2 1198 1 1195
2 1199 1 1195
2 1201 1 1200
2 1202 1 1200
2 1203 1 1200
2 1204 1 1200
2 1206 1 1205
2 1207 1 1205
2 1208 1 1205
2 1209 1 1205
2 1217 1 1216
2 1218 1 1216
2 1220 1 1219
2 1221 1 1219
2 1223 1 1222
2 1224 1 1222
2 1226 1 1225
2 1227 1 1225
2 1229 1 1228
2 1230 1 1228
2 1232 1 1231
2 1233 1 1231
2 1235 1 1234
2 1236 1 1234
2 1238 1 1237
2 1239 1 1237
2 1241 1 1240
2 1242 1 1240
2 1244 1 1243
2 1245 1 1243
2 1247 1 1246
2 1248 1 1246
2 1252 1 1251
2 1253 1 1251
2 1255 1 1254
2 1256 1 1254
2 1258 1 1257
2 1259 1 1257
2 1261 1 1260
2 1262 1 1260
2 1264 1 1263
2 1265 1 1263
2 1267 1 1266
2 1268 1 1266
2 1497 1 1496
2 1498 1 1496
2 1500 1 1499
2 1501 1 1499
2 1503 1 1502
2 1504 1 1502
2 1505 1 1502
2 1507 1 1506
2 1508 1 1506
2 1509 1 1506
2 1511 1 1510
2 1512 1 1510
2 1514 1 1513
2 1515 1 1513
2 1517 1 1516
2 1518 1 1516
2 1554 1 1553
2 1555 1 1553
2 1556 1 1553
2 1558 1 1557
2 1559 1 1557
2 1560 1 1557
2 1562 1 1561
2 1563 1 1561
2 1579 1 1578
2 1580 1 1578
2 1583 1 1582
2 1584 1 1582
2 1586 1 1585
2 1587 1 1585
2 1589 1 1588
2 1590 1 1588
2 1592 1 1591
2 1593 1 1591
2 1594 1 1591
2 1595 1 1591
2 1597 1 1596
2 1598 1 1596
2 1599 1 1596
2 1601 1 1600
2 1602 1 1600
2 1603 1 1600
2 1604 1 1600
2 1605 1 1600
2 1607 1 1606
2 1608 1 1606
2 1609 1 1606
2 1610 1 1606
2 1611 1 1606
2 1613 1 1612
2 1614 1 1612
2 1616 1 1615
2 1617 1 1615
2 1618 1 1615
2 1620 1 1619
2 1621 1 1619
2 1622 1 1619
2 1623 1 1619
2 1625 1 1624
2 1626 1 1624
2 1627 1 1624
2 1629 1 1628
2 1630 1 1628
2 1632 1 1631
2 1633 1 1631
2 1635 1 1634
2 1636 1 1634
2 1638 1 1637
2 1639 1 1637
2 1640 1 1637
2 1641 1 1637
2 1643 1 1642
2 1644 1 1642
2 1645 1 1642
2 1646 1 1642
2 1648 1 1647
2 1649 1 1647
2 1650 1 1647
2 1652 1 1651
2 1653 1 1651
2 1654 1 1651
2 1655 1 1651
2 1657 1 1656
2 1658 1 1656
2 1659 1 1656
2 1677 1 1676
2 1678 1 1676
2 1679 1 1676
2 1680 1 1676
2 1682 1 1681
2 1683 1 1681
2 1684 1 1681
2 1685 1 1681
2 1687 1 1686
2 1688 1 1686
2 1689 1 1686
2 1691 1 1690
2 1692 1 1690
2 1709 1 1708
2 1710 1 1708
2 1771 1 1770
2 1772 1 1770
2 1774 1 1773
2 1775 1 1773
2 1779 1 1778
2 1780 1 1778
2 1782 1 1781
2 1783 1 1781
2 1796 1 1795
2 1797 1 1795
2 1799 1 1798
2 1800 1 1798
2 1802 1 1801
2 1803 1 1801
2 1805 1 1804
2 1806 1 1804
2 1825 1 1824
2 1826 1 1824
2 1828 1 1827
2 1829 1 1827
2 1834 1 1833
2 1835 1 1833
2 1837 1 1836
2 1838 1 1836
2 1839 1 1836
2 1840 1 1836
2 1842 1 1841
2 1843 1 1841
2 1844 1 1841
2 1845 1 1841
2 1846 1 1841
2 1847 1 1841
2 1849 1 1848
2 1850 1 1848
2 1851 1 1848
2 1853 1 1852
2 1854 1 1852
2 1855 1 1852
2 1857 1 1856
2 1858 1 1856
2 1859 1 1856
2 1860 1 1856
2 1861 1 1856
2 1862 1 1856
2 1864 1 1863
2 1865 1 1863
2 1866 1 1863
2 1867 1 1863
2 1868 1 1863
2 1869 1 1863
2 1871 1 1870
2 1872 1 1870
2 1873 1 1870
2 1874 1 1870
2 1876 1 1875
2 1877 1 1875
2 1878 1 1875
2 1879 1 1875
2 1881 1 1880
2 1882 1 1880
2 1883 1 1880
2 1884 1 1880
2 1886 1 1885
2 1887 1 1885
2 1889 1 1888
2 1890 1 1888
2 1892 1 1891
2 1893 1 1891
2 1895 1 1894
2 1896 1 1894
2 1898 1 1897
2 1899 1 1897
2 1937 1 1936
2 1938 1 1936
2 1943 1 1942
2 1944 1 1942
2 1946 1 1945
2 1947 1 1945
2 1949 1 1948
2 1950 1 1948
2 1952 1 1951
2 1953 1 1951
2 1955 1 1954
2 1956 1 1954
2 1958 1 1957
2 1959 1 1957
2 1961 1 1960
2 1962 1 1960
2 1964 1 1963
2 1965 1 1963
2 1967 1 1966
2 1968 1 1966
2 2047 1 2046
2 2048 1 2046
2 2050 1 2049
2 2051 1 2049
2 2053 1 2052
2 2054 1 2052
2 2056 1 2055
2 2057 1 2055
2 2059 1 2058
2 2060 1 2058
2 2062 1 2061
2 2063 1 2061
2 2065 1 2064
2 2066 1 2064
2 2068 1 2067
2 2069 1 2067
2 2071 1 2070
2 2072 1 2070
2 2074 1 2073
2 2075 1 2073
2 2077 1 2076
2 2078 1 2076
2 2080 1 2079
2 2081 1 2079
2 2096 1 2095
2 2097 1 2095
2 2099 1 2098
2 2100 1 2098
2 2102 1 2101
2 2103 1 2101
2 2105 1 2104
2 2106 1 2104
2 2108 1 2107
2 2109 1 2107
2 2111 1 2110
2 2112 1 2110
2 2114 1 2113
2 2115 1 2113
2 2116 1 2113
2 2117 1 2113
2 2118 1 2113
2 2121 1 2120
2 2122 1 2120
2 2123 1 2120
2 2124 1 2120
2 2129 1 2128
2 2130 1 2128
2 2131 1 2128
2 2132 1 2128
2 2133 1 2128
2 2134 1 2128
2 2136 1 2135
2 2137 1 2135
2 2138 1 2135
2 2139 1 2135
2 2140 1 2135
2 2142 1 2141
2 2143 1 2141
2 2145 1 2144
2 2146 1 2144
2 2148 1 2147
2 2149 1 2147
2 2151 1 2150
2 2152 1 2150
2 2186 1 2185
2 2187 1 2185
2 2189 1 2188
2 2190 1 2188
2 2192 1 2191
2 2193 1 2191
2 2195 1 2194
2 2196 1 2194
2 2198 1 2197
2 2199 1 2197
2 2202 1 2201
2 2203 1 2201
2 2205 1 2204
2 2206 1 2204
2 2208 1 2207
2 2209 1 2207
2 2211 1 2210
2 2212 1 2210
2 2214 1 2213
2 2215 1 2213
2 2217 1 2216
2 2218 1 2216
2 2220 1 2219
2 2221 1 2219
2 2251 1 2250
2 2252 1 2250
2 2267 1 2266
2 2268 1 2266
2 2270 1 2269
2 2271 1 2269
2 2292 1 2291
2 2293 1 2291
2 2295 1 2294
2 2296 1 2294
2 2360 1 2359
2 2361 1 2359
2 2369 1 2368
2 2370 1 2368
2 2371 1 2368
2 2378 1 2377
2 2379 1 2377
2 2380 1 2377
2 2381 1 2377
2 2383 1 2382
2 2384 1 2382
2 2385 1 2382
2 2392 1 2391
2 2393 1 2391
2 2394 1 2391
2 2396 1 2395
2 2397 1 2395
2 2398 1 2395
2 2399 1 2395
2 2418 1 2417
2 2419 1 2417
2 2420 1 2417
2 2422 1 2421
2 2423 1 2421
2 2424 1 2421
2 2426 1 2425
2 2427 1 2425
2 2435 1 2434
2 2436 1 2434
2 2438 1 2437
2 2439 1 2437
2 2441 1 2440
2 2442 1 2440
2 2444 1 2443
2 2445 1 2443
2 2447 1 2446
2 2448 1 2446
2 2450 1 2449
2 2451 1 2449
2 2455 1 2454
2 2456 1 2454
2 2458 1 2457
2 2459 1 2457
2 2461 1 2460
2 2462 1 2460
2 2464 1 2463
2 2465 1 2463
2 2467 1 2466
2 2468 1 2466
2 2470 1 2469
2 2471 1 2469
2 2473 1 2472
2 2474 1 2472
2 2476 1 2475
2 2477 1 2475
2 2479 1 2478
2 2480 1 2478
2 2482 1 2481
2 2483 1 2481
2 2485 1 2484
2 2486 1 2484
2 2488 1 2487
2 2489 1 2487
2 2491 1 2490
2 2492 1 2490
2 2494 1 2493
2 2495 1 2493
2 2522 1 2521
2 2523 1 2521
2 2532 1 2531
2 2533 1 2531
2 2535 1 2534
2 2536 1 2534
2 2538 1 2537
2 2539 1 2537
2 2541 1 2540
2 2542 1 2540
2 2604 1 2603
2 2605 1 2603
2 2606 1 2603
2 2614 1 2613
2 2615 1 2613
2 2616 1 2613
2 2622 1 2621
2 2623 1 2621
2 2625 1 2624
2 2626 1 2624
2 2627 1 2624
2 2639 1 2638
2 2640 1 2638
2 2641 1 2638
2 2642 1 2638
2 2647 1 2646
2 2648 1 2646
2 2649 1 2646
2 2650 1 2646
2 2660 1 2659
2 2661 1 2659
2 2662 1 2659
2 2682 1 2681
2 2683 1 2681
2 2685 1 2684
2 2686 1 2684
2 2688 1 2687
2 2689 1 2687
2 2691 1 2690
2 2692 1 2690
2 2704 1 2703
2 2705 1 2703
2 2730 1 2729
2 2731 1 2729
2 2732 1 2729
2 2733 1 2729
2 2739 1 2738
2 2740 1 2738
2 2741 1 2738
2 2742 1 2738
2 2762 1 2761
2 2763 1 2761
2 2764 1 2761
2 2765 1 2761
2 2767 1 2766
2 2768 1 2766
2 2769 1 2766
2 2770 1 2766
2 2794 1 2793
2 2795 1 2793
2 2797 1 2796
2 2798 1 2796
2 2799 1 2796
2 2801 1 2800
2 2802 1 2800
2 2804 1 2803
2 2805 1 2803
2 2807 1 2806
2 2808 1 2806
2 2818 1 2817
2 2819 1 2817
2 2821 1 2820
2 2822 1 2820
2 2823 1 2820
2 2824 1 2820
2 2825 1 2820
2 2827 1 2826
2 2828 1 2826
2 2832 1 2831
2 2833 1 2831
2 2834 1 2831
2 2835 1 2831
2 2836 1 2831
2 2842 1 2841
2 2843 1 2841
2 2845 1 2844
2 2846 1 2844
2 2847 1 2844
2 2848 1 2844
2 2849 1 2844
2 2855 1 2854
2 2856 1 2854
2 2857 1 2854
2 2858 1 2854
2 2860 1 2859
2 2861 1 2859
2 2862 1 2859
2 2863 1 2859
2 2864 1 2859
2 2870 1 2869
2 2871 1 2869
2 2872 1 2869
2 2873 1 2869
2 2875 1 2874
2 2876 1 2874
2 2878 1 2877
2 2879 1 2877
2 2883 1 2882
2 2884 1 2882
2 2886 1 2885
2 2887 1 2885
2 2889 1 2888
2 2890 1 2888
2 2932 1 2931
2 2933 1 2931
2 2973 1 2972
2 2974 1 2972
2 2976 1 2975
2 2977 1 2975
2 2979 1 2978
2 2980 1 2978
2 2982 1 2981
2 2983 1 2981
2 2987 1 2986
2 2988 1 2986
2 2990 1 2989
2 2991 1 2989
2 2993 1 2992
2 2994 1 2992
2 2996 1 2995
2 2997 1 2995
2 2999 1 2998
2 3000 1 2998
2 3002 1 3001
2 3003 1 3001
2 3005 1 3004
2 3006 1 3004
2 3011 1 3010
2 3012 1 3010
2 3014 1 3013
2 3015 1 3013
2 3017 1 3016
2 3018 1 3016
2 3020 1 3019
2 3021 1 3019
2 3023 1 3022
2 3024 1 3022
2 3026 1 3025
2 3027 1 3025
2 3031 1 3030
2 3032 1 3030
2 3033 1 3030
2 3034 1 3030
2 3040 1 3039
2 3041 1 3039
2 3042 1 3039
2 3043 1 3039
2 3051 1 3050
2 3052 1 3050
2 3062 1 3061
2 3063 1 3061
2 3077 1 3076
2 3078 1 3076
2 3089 1 3088
2 3090 1 3088
2 3092 1 3091
2 3093 1 3091
2 3111 1 3110
2 3112 1 3110
2 3114 1 3113
2 3115 1 3113
2 3138 1 3137
2 3139 1 3137
2 3141 1 3140
2 3142 1 3140
2 3144 1 3143
2 3145 1 3143
2 3147 1 3146
2 3148 1 3146
2 3150 1 3149
2 3151 1 3149
2 3153 1 3152
2 3154 1 3152
2 3158 1 3157
2 3159 1 3157
2 3161 1 3160
2 3162 1 3160
2 3164 1 3163
2 3165 1 3163
2 3167 1 3166
2 3168 1 3166
2 3170 1 3169
2 3171 1 3169
2 3173 1 3172
2 3174 1 3172
2 3181 1 3180
2 3182 1 3180
2 3239 1 3238
2 3240 1 3238
2 3242 1 3241
2 3243 1 3241
2 3245 1 3244
2 3246 1 3244
2 3248 1 3247
2 3249 1 3247
2 3251 1 3250
2 3252 1 3250
2 3254 1 3253
2 3255 1 3253
2 3257 1 3256
2 3258 1 3256
2 3260 1 3259
2 3261 1 3259
2 3263 1 3262
2 3264 1 3262
2 3266 1 3265
2 3267 1 3265
2 3269 1 3268
2 3270 1 3268
2 3272 1 3271
2 3273 1 3271
2 3275 1 3274
2 3276 1 3274
2 3278 1 3277
2 3279 1 3277
2 3316 1 3315
2 3317 1 3315
2 3319 1 3318
2 3320 1 3318
2 3322 1 3321
2 3323 1 3321
2 3325 1 3324
2 3326 1 3324
2 3328 1 3327
2 3329 1 3327
2 3331 1 3330
2 3332 1 3330
2 3341 1 3340
2 3342 1 3340
2 3345 1 3344
2 3346 1 3344
2 3349 1 3348
2 3350 1 3348
2 3353 1 3352
2 3354 1 3352
2 3357 1 3356
2 3358 1 3356
2 3361 1 3360
2 3362 1 3360
2 3365 1 3364
2 3366 1 3364
2 3368 1 3367
2 3369 1 3367
2 3371 1 3370
2 3372 1 3370
2 3375 1 3374
2 3376 1 3374
2 3379 1 3378
2 3380 1 3378
2 3383 1 3382
2 3384 1 3382
2 3387 1 3386
2 3388 1 3386
2 3391 1 3390
2 3392 1 3390
2 3395 1 3394
2 3396 1 3394
2 3398 1 3397
2 3399 1 3397
2 3451 1 3450
2 3452 1 3450
2 3454 1 3453
2 3455 1 3453
2 3457 1 3456
2 3458 1 3456
2 3460 1 3459
2 3461 1 3459
2 3523 1 3522
2 3524 1 3522
2 3526 1 3525
2 3527 1 3525
2 3529 1 3528
2 3530 1 3528
2 3532 1 3531
2 3533 1 3531
2 3535 1 3534
2 3536 1 3534
2 3538 1 3537
2 3539 1 3537
2 3541 1 3540
2 3542 1 3540
2 3544 1 3543
2 3545 1 3543
2 3577 1 3576
2 3578 1 3576
2 3580 1 3579
2 3581 1 3579
2 3586 1 3585
2 3587 1 3585
2 3589 1 3588
2 3590 1 3588
2 3601 1 3600
2 3602 1 3600
2 3604 1 3603
2 3605 1 3603
2 3606 1 3603
2 3607 1 3603
2 3609 1 3608
2 3610 1 3608
2 3611 1 3608
2 3613 1 3612
2 3614 1 3612
2 3617 1 3616
2 3618 1 3616
2 3619 1 3616
2 3620 1 3616
2 3621 1 3616
2 3623 1 3622
2 3624 1 3622
2 3625 1 3622
2 3626 1 3622
2 3636 1 3635
2 3637 1 3635
2 3638 1 3635
2 3639 1 3635
2 3641 1 3640
2 3642 1 3640
2 3643 1 3640
2 3645 1 3644
2 3646 1 3644
2 3649 1 3648
2 3650 1 3648
2 3651 1 3648
2 3652 1 3648
2 3653 1 3648
2 3655 1 3654
2 3656 1 3654
2 3657 1 3654
2 3658 1 3654
2 3724 1 3723
2 3725 1 3723
2 3738 1 3737
2 3739 1 3737
2 3755 1 3754
2 3756 1 3754
2 3757 1 3754
2 3759 1 3758
2 3760 1 3758
2 3763 1 3762
2 3764 1 3762
2 3768 1 3767
2 3769 1 3767
2 3770 1 3767
2 3772 1 3771
2 3773 1 3771
2 3776 1 3775
2 3777 1 3775
2 3781 1 3780
2 3782 1 3780
2 3791 1 3790
2 3792 1 3790
2 3824 1 3823
2 3825 1 3823
2 3828 1 3827
2 3829 1 3827
2 3841 1 3840
2 3842 1 3840
2 3844 1 3843
2 3845 1 3843
2 3846 1 3843
2 3853 1 3852
2 3854 1 3852
2 3860 1 3859
2 3861 1 3859
2 3865 1 3864
2 3866 1 3864
2 3871 1 3870
2 3872 1 3870
2 3878 1 3877
2 3879 1 3877
