1 1 0 2 0
1 4 0 6 0
1 11 0 2 0
1 14 0 2 0
1 17 0 2 0
1 20 0 2 0
1 23 0 1 0
1 24 0 1 0
1 25 0 1 0
1 26 0 1 0
1 27 0 3 0
1 31 0 2 0
1 34 0 2 0
1 37 0 2 0
1 40 0 2 0
1 43 0 2 0
1 46 0 2 0
1 49 0 2 0
1 52 0 1 0
1 53 0 1 0
1 54 0 6 0
1 61 0 2 0
1 64 0 2 0
1 67 0 2 0
1 70 0 2 0
1 73 0 2 0
1 76 0 2 0
1 79 0 1 0
1 80 0 1 0
1 81 0 1 0
1 82 0 1 0
1 83 0 2 0
1 86 0 1 0
1 87 0 1 0
1 88 0 2 0
1 91 0 2 0
1 94 0 2 0
1 97 0 2 0
1 100 0 2 0
1 103 0 2 0
1 106 0 2 0
1 109 0 2 0
1 112 0 1 0
1 113 0 1 0
1 114 0 1 0
1 115 0 1 0
1 116 0 1 0
1 117 0 1 0
1 118 0 1 0
1 119 0 1 0
1 120 0 1 0
1 121 0 1 0
1 122 0 1 0
1 123 0 2 0
1 126 0 1 0
1 127 0 1 0
1 128 0 1 0
1 129 0 1 0
1 130 0 1 0
1 131 0 1 0
1 132 0 2 0
1 135 0 1 0
1 136 0 1 0
1 137 0 2 0
1 140 0 1 0
1 141 0 3 0
1 145 0 1 0
1 146 0 2 0
1 149 0 2 0
1 152 0 2 0
1 155 0 2 0
1 158 0 2 0
1 161 0 2 0
1 164 0 2 0
1 167 0 2 0
1 170 0 2 0
1 173 0 2 0
1 176 0 2 0
1 179 0 2 0
1 182 0 2 0
1 185 0 2 0
1 188 0 2 0
1 191 0 2 0
1 194 0 2 0
1 197 0 2 0
1 200 0 2 0
1 203 0 2 0
1 206 0 2 0
1 209 0 1 0
1 210 0 6 0
1 217 0 1 0
1 218 0 6 0
1 225 0 1 0
1 226 0 6 0
1 233 0 1 0
1 234 0 6 0
1 241 0 1 0
1 242 0 2 0
1 245 0 2 0
1 248 0 2 0
1 251 0 2 0
1 254 0 2 0
1 257 0 6 0
1 264 0 1 0
1 265 0 6 0
1 272 0 1 0
1 273 0 6 0
1 280 0 1 0
1 281 0 6 0
1 288 0 1 0
1 289 0 2 0
1 292 0 1 0
1 293 0 5 0
1 299 0 2 0
1 302 0 4 0
1 307 0 1 0
1 308 0 6 0
1 315 0 1 0
1 316 0 6 0
1 323 0 1 0
1 324 0 6 0
1 331 0 1 0
1 332 0 2 0
1 335 0 2 0
1 338 0 2 0
1 341 0 6 0
1 348 0 2 0
1 351 0 6 0
1 358 0 2 0
1 361 0 4 0
1 366 0 2 0
1 369 0 2 0
1 372 0 1 0
1 373 0 1 0
1 374 0 11 0
1 386 0 2 0
1 389 0 10 0
1 400 0 10 0
1 411 0 10 0
1 422 0 12 0
1 435 0 10 0
1 446 0 10 0
1 457 0 10 0
1 468 0 10 0
1 479 0 10 0
1 490 0 12 0
1 503 0 10 0
1 514 0 8 0
1 523 0 10 0
1 534 0 10 0
1 545 0 3 0
1 549 0 2 0
1 552 0 3 0
1 556 0 2 0
1 559 0 2 0
1 562 0 3 0
1 566 0 4 0
1 571 0 2 0
1 574 0 2 0
1 577 0 2 0
1 580 0 2 0
1 583 0 4 0
1 588 0 2 0
1 591 0 1 0
1 592 0 2 0
1 595 0 1 0
1 596 0 1 0
1 597 0 1 0
1 598 0 1 0
1 599 0 3 0
1 603 0 3 0
1 607 0 2 0
1 610 0 2 0
1 613 0 2 0
1 616 0 2 0
1 619 0 5 0
1 625 0 5 0
1 631 0 1 0
3 709 9 0 1 142
3 816 9 0 1 294
0 1042 7 1 2 135 631
0 1043 5 1 1 591
3 1066 9 0 1 593
0 1067 5 12 1 595
0 1080 5 11 1 596
0 1092 5 11 1 597
0 1104 5 12 1 598
3 1137 5 0 1 546
3 1138 5 0 1 349
3 1139 5 0 1 367
3 1140 7 0 2 553 563
3 1141 5 0 1 550
3 1142 5 0 1 547
3 1143 5 0 1 548
3 1144 5 0 1 339
3 1145 5 0 1 359
0 1146 6 1 2 373 2
3 1147 7 0 2 143 145
0 1148 5 1 1 594
0 1149 5 1 1 1042
0 1150 7 1 2 1043 28
0 1151 7 1 2 387 557
3 1152 5 0 1 246
3 1153 5 0 1 554
3 1154 5 0 1 564
3 1155 5 0 1 560
0 1156 7 1 4 388 561 558 555
0 1157 5 3 1 567
0 1161 9 11 1 572
0 1173 9 11 1 575
0 1185 9 11 1 573
0 1197 9 11 1 576
0 1209 9 3 1 138
0 1213 9 2 1 139
0 1216 9 2 1 144
0 1219 5 3 1 584
0 1223 9 11 1 578
0 1235 9 11 1 581
0 1247 9 11 1 579
0 1259 9 11 1 582
0 1271 9 8 1 255
0 1280 9 11 1 252
0 1292 9 10 1 253
0 1303 9 11 1 249
0 1315 9 11 1 250
0 1327 9 11 1 611
0 1339 9 11 1 608
0 1351 9 11 1 614
0 1363 9 11 1 617
0 1375 9 2 1 211
0 1378 9 2 1 212
0 1381 9 2 1 219
0 1384 9 2 1 220
0 1387 9 2 1 227
0 1390 9 2 1 228
0 1393 9 2 1 235
0 1396 9 2 1 236
0 1415 9 2 1 258
0 1418 9 2 1 259
0 1421 9 2 1 266
0 1424 9 2 1 267
0 1427 9 2 1 274
0 1430 9 2 1 275
0 1433 9 2 1 282
0 1436 9 2 1 283
0 1455 9 6 1 336
0 1462 9 6 1 337
0 1469 9 5 1 207
0 1475 7 3 2 29 32
0 1479 9 2 1 3
0 1482 9 9 1 589
0 1492 9 2 1 295
0 1495 9 2 1 303
0 1498 9 2 1 309
0 1501 9 2 1 310
0 1504 9 2 1 317
0 1507 9 2 1 318
0 1510 9 2 1 325
0 1513 9 2 1 326
0 1516 9 2 1 342
0 1519 9 2 1 343
0 1522 9 2 1 352
0 1525 9 2 1 353
0 1542 9 2 1 260
0 1545 9 2 1 261
0 1548 9 2 1 268
0 1551 9 2 1 269
0 1554 9 2 1 276
0 1557 9 2 1 277
0 1560 9 2 1 284
0 1563 9 2 1 285
0 1566 9 6 1 333
0 1573 9 6 1 334
0 1580 9 2 1 551
0 1583 7 4 2 33 30
0 1588 5 5 1 590
0 1594 9 2 1 327
0 1597 9 2 1 328
0 1600 9 2 1 344
0 1603 9 2 1 345
0 1606 9 2 1 354
0 1609 9 2 1 355
0 1612 9 2 1 296
0 1615 9 2 1 304
0 1618 9 2 1 311
0 1621 9 2 1 312
0 1624 9 2 1 319
0 1627 9 2 1 320
0 1630 9 2 1 362
0 1633 9 2 1 363
0 1636 9 2 1 213
0 1639 9 2 1 214
0 1642 9 2 1 221
0 1645 9 2 1 222
0 1648 9 2 1 229
0 1651 9 2 1 230
0 1654 9 2 1 237
0 1657 9 2 1 238
0 1660 5 2 1 329
0 1663 9 11 1 243
0 1675 9 9 1 244
0 1685 9 11 1 256
0 1697 9 11 1 612
0 1709 9 11 1 609
0 1721 9 5 1 626
0 1727 9 3 1 620
0 1731 9 11 1 615
0 1743 9 11 1 618
0 1755 5 2 1 600
0 1758 5 2 1 604
0 1761 9 7 1 621
0 1769 9 7 1 627
0 1777 9 7 1 622
0 1785 9 7 1 628
0 1793 9 6 1 623
0 1800 9 6 1 629
0 1807 9 6 1 624
0 1814 9 6 1 630
0 1821 9 2 1 300
0 1824 9 2 1 447
0 1827 9 2 1 458
0 1830 9 2 1 469
0 1833 9 2 1 423
0 1836 9 2 1 436
0 1839 9 2 1 390
0 1842 9 2 1 401
0 1845 9 2 1 412
0 1848 9 2 1 375
0 1851 9 2 1 5
0 1854 9 2 1 448
0 1857 9 2 1 459
0 1860 9 2 1 470
0 1863 9 2 1 437
0 1866 9 2 1 391
0 1869 9 2 1 402
0 1872 9 2 1 413
0 1875 9 2 1 424
0 1878 9 2 1 376
0 1881 9 2 1 480
0 1884 9 2 1 491
0 1887 9 2 1 504
0 1890 9 2 1 515
0 1893 9 2 1 524
0 1896 9 2 1 535
0 1899 9 2 1 55
0 1902 9 2 1 481
0 1905 9 2 1 505
0 1908 9 2 1 516
0 1911 9 2 1 525
0 1914 9 2 1 536
0 1917 9 2 1 492
0 1920 9 2 1 364
0 1923 9 2 1 370
0 1926 9 2 1 346
0 1929 9 2 1 356
0 1932 9 2 1 313
0 1935 9 2 1 321
0 1938 9 2 1 297
0 1941 9 2 1 305
0 1944 9 2 1 286
0 1947 9 2 1 290
0 1950 9 2 1 270
0 1953 9 2 1 278
0 1956 9 2 1 239
0 1959 9 2 1 262
0 1962 9 2 1 223
0 1965 9 2 1 231
0 1968 9 2 1 215
3 1972 5 0 1 1146
3 2054 7 0 2 136 1148
3 2060 5 0 1 1150
3 2061 5 0 1 1151
3 2139 9 0 1 1210
3 2142 9 0 1 1217
3 2309 9 0 1 1480
0 2349 7 1 2 1105 517
0 2350 3 1 2 1068 518
3 2387 9 0 1 1581
3 2527 9 0 1 1822
3 2584 5 0 1 1582
0 2585 7 1 3 171 1162 1174
0 2586 7 1 3 174 1163 1175
0 2587 7 1 3 168 1164 1176
0 2588 7 1 3 165 1165 1177
0 2589 7 1 3 162 1166 1178
3 2590 6 0 2 1476 140
0 2591 7 1 3 186 1186 1198
0 2592 7 1 3 159 1187 1199
0 2593 7 1 3 153 1188 1200
0 2594 7 1 3 147 1189 1201
0 2595 7 1 3 172 1224 1236
0 2596 7 1 3 175 1225 1237
0 2597 7 1 3 169 1226 1238
0 2598 7 1 3 166 1227 1239
0 2599 7 1 3 163 1228 1240
0 2600 7 1 3 187 1248 1260
0 2601 7 1 3 160 1249 1261
0 2602 7 1 3 154 1250 1262
0 2603 7 1 3 148 1251 1263
0 2604 7 1 3 107 1732 1744
0 2605 7 1 3 62 1328 1340
0 2606 7 1 3 108 1698 1710
0 2607 7 1 3 50 1699 1711
0 2608 7 1 3 104 1700 1712
0 2609 7 1 3 41 1701 1713
0 2610 7 1 3 38 1702 1714
0 2611 7 1 3 21 1329 1341
0 2612 7 1 3 18 1330 1342
0 2613 7 1 3 71 1331 1343
0 2614 7 1 3 65 1332 1344
0 2615 7 1 3 51 1733 1745
0 2616 7 1 3 105 1734 1746
0 2617 7 1 3 42 1735 1747
0 2618 7 1 3 39 1736 1748
0 2619 7 1 3 22 1352 1364
0 2620 7 1 3 19 1353 1365
0 2621 7 1 3 72 1354 1366
0 2622 7 1 3 66 1355 1367
3 2623 5 0 1 1477
0 2624 7 1 3 124 1759 601
0 2625 7 1 2 1778 1786
0 2626 7 1 3 63 1356 1368
0 2627 7 1 2 1762 1770
0 2628 5 1 1 1825
0 2629 5 1 1 1828
0 2630 5 1 1 1831
0 2631 5 1 1 1834
0 2632 5 1 1 1837
0 2633 5 1 1 1840
0 2634 5 1 1 1843
0 2635 5 1 1 1846
0 2636 5 1 1 1849
0 2637 5 1 1 1852
0 2638 5 1 1 1855
0 2639 5 1 1 1858
0 2640 5 1 1 1861
0 2641 5 1 1 1864
0 2642 5 1 1 1867
0 2643 5 1 1 1870
0 2644 5 1 1 1873
0 2645 5 1 1 1876
0 2646 5 1 1 1879
0 2647 9 5 1 1211
0 2653 5 10 1 1167
0 2664 5 10 1 1179
0 2675 9 5 1 1212
0 2681 5 10 1 1190
0 2692 5 10 1 1202
0 2703 7 1 3 180 1191 1203
0 2704 9 4 1 1481
0 2709 5 1 1 1882
0 2710 5 1 1 1885
0 2711 5 1 1 1888
0 2712 5 1 1 1891
0 2713 5 1 1 1894
0 2714 5 1 1 1897
0 2715 5 1 1 1900
0 2716 5 1 1 1903
0 2717 5 1 1 1906
0 2718 5 1 1 1909
0 2719 5 1 1 1912
0 2720 5 1 1 1915
0 2721 5 1 1 1918
0 2722 9 5 1 1214
0 2728 5 10 1 1229
0 2739 5 10 1 1241
0 2750 9 5 1 1215
0 2756 5 10 1 1252
0 2767 5 10 1 1264
0 2778 7 1 3 181 1253 1265
0 2779 5 10 1 1333
0 2790 5 10 1 1345
0 2801 5 10 1 1357
0 2812 5 10 1 1369
0 2823 5 1 1 1376
0 2824 5 1 1 1379
0 2825 5 1 1 1382
0 2826 5 1 1 1385
0 2827 5 1 1 1388
0 2828 5 1 1 1391
0 2829 5 1 1 1394
0 2830 5 1 1 1397
0 2831 7 1 3 1106 460 1380
0 2832 7 1 3 1107 471 1386
0 2833 7 1 3 1108 425 1392
0 2834 7 1 3 1109 438 1398
0 2835 7 1 2 1069 1377
0 2836 7 1 2 1070 1383
0 2837 7 1 2 1071 1389
0 2838 7 1 2 1072 1395
0 2839 5 1 1 1416
0 2840 5 1 1 1419
0 2841 5 1 1 1422
0 2842 5 1 1 1425
0 2843 5 1 1 1428
0 2844 5 1 1 1431
0 2845 5 1 1 1434
0 2846 5 1 1 1437
0 2847 7 1 3 1110 392 1420
0 2848 7 1 3 1111 403 1426
0 2849 7 1 3 1112 414 1432
0 2850 7 1 3 1113 377 1438
0 2851 7 1 2 1073 1417
0 2852 7 1 2 1074 1423
0 2853 7 1 2 1075 1429
0 2854 7 1 2 1076 1435
0 2855 5 5 1 1456
0 2861 5 5 1 1463
0 2867 7 1 2 292 1457
0 2868 7 1 2 288 1458
0 2869 7 1 2 280 1459
0 2870 7 1 2 272 1460
0 2871 7 1 2 264 1461
0 2872 7 1 2 241 1464
0 2873 7 1 2 233 1465
0 2874 7 1 2 225 1466
0 2875 7 1 2 217 1467
0 2876 7 1 2 209 1468
0 2877 9 4 1 1218
0 2882 5 8 1 1483
0 2891 5 9 1 1478
0 2901 5 1 1 1493
0 2902 5 1 1 1496
0 2903 5 1 1 1499
0 2904 5 1 1 1502
0 2905 5 1 1 1505
0 2906 5 1 1 1508
0 2907 7 1 2 1304 1497
0 2908 7 1 3 1305 482 1503
0 2909 7 1 3 1306 493 1509
0 2910 7 1 2 1664 1494
0 2911 7 1 2 1665 1500
0 2912 7 1 2 1666 1506
0 2913 5 1 1 1511
0 2914 5 1 1 1514
0 2915 5 1 1 1517
0 2916 5 1 1 1520
0 2917 5 1 1 1523
0 2918 5 1 1 1526
0 2919 7 1 3 1114 506 1515
0 2920 5 1 1 2349
0 2921 7 1 3 1115 526 1521
0 2922 7 1 3 1116 537 1527
0 2923 7 1 2 1077 1512
0 2924 7 1 2 1078 1518
0 2925 7 1 2 1079 1524
0 2926 5 1 1 1543
0 2927 5 1 1 1546
0 2928 5 1 1 1549
0 2929 5 1 1 1552
0 2930 5 1 1 1555
0 2931 5 1 1 1558
0 2932 5 1 1 1561
0 2933 5 1 1 1564
0 2934 7 1 3 1307 393 1547
0 2935 7 1 3 1308 404 1553
0 2936 7 1 3 1309 415 1559
0 2937 7 1 3 1310 378 1565
0 2938 7 1 2 1667 1544
0 2939 7 1 2 1668 1550
0 2940 7 1 2 1669 1556
0 2941 7 1 2 1670 1562
0 2942 5 5 1 1567
0 2948 5 5 1 1574
0 2954 7 1 2 372 1568
0 2955 7 1 2 368 1569
0 2956 7 1 2 360 1570
0 2957 7 1 2 350 1571
0 2958 7 1 2 340 1572
0 2959 7 1 2 331 1575
0 2960 7 1 2 323 1576
0 2961 7 1 2 315 1577
0 2962 7 1 2 307 1578
0 2963 7 1 2 301 1579
0 2964 5 4 1 1589
0 2969 7 1 2 84 1590
0 2970 7 1 2 86 1591
0 2971 7 1 2 89 1592
0 2972 7 1 2 90 1593
0 2973 5 1 1 1595
0 2974 5 1 1 1598
0 2975 5 1 1 1601
0 2976 5 1 1 1604
0 2977 5 1 1 1607
0 2978 5 1 1 1610
0 2979 7 1 3 1316 507 1599
0 2980 7 1 2 1317 519
0 2981 7 1 3 1318 527 1605
0 2982 7 1 3 1319 538 1611
0 2983 7 1 2 1676 1596
0 2984 3 1 2 1677 520
0 2985 7 1 2 1678 1602
0 2986 7 1 2 1679 1608
0 2987 5 1 1 1613
0 2988 5 1 1 1616
0 2989 5 1 1 1619
0 2990 5 1 1 1622
0 2991 5 1 1 1625
0 2992 5 1 1 1628
0 2993 7 1 2 1320 1617
0 2994 7 1 3 1321 483 1623
0 2995 7 1 3 1322 494 1629
0 2996 7 1 2 1680 1614
0 2997 7 1 2 1681 1620
0 2998 7 1 2 1682 1626
0 2999 5 1 1 1631
0 3000 9 2 1 1470
0 3003 9 2 1 1471
0 3006 5 1 1 1634
0 3007 9 2 1 1472
0 3010 9 2 1 1473
0 3013 7 1 2 1323 1632
0 3014 7 1 2 1324 1635
0 3015 5 1 1 1637
0 3016 5 1 1 1640
0 3017 5 1 1 1643
0 3018 5 1 1 1646
0 3019 5 1 1 1649
0 3020 5 1 1 1652
0 3021 5 1 1 1655
0 3022 5 1 1 1658
0 3023 7 1 3 1311 461 1641
0 3024 7 1 3 1312 472 1647
0 3025 7 1 3 1313 426 1653
0 3026 7 1 3 1314 439 1659
0 3027 7 1 2 1671 1638
0 3028 7 1 2 1672 1644
0 3029 7 1 2 1673 1650
0 3030 7 1 2 1674 1656
0 3031 5 1 1 1921
0 3032 5 1 1 1924
0 3033 5 1 1 1927
0 3034 5 1 1 1930
0 3035 9 2 1 1661
0 3038 9 2 1 1662
0 3041 5 10 1 1703
0 3052 5 10 1 1715
0 3063 5 4 1 1722
0 3068 5 2 1 1728
0 3071 7 1 2 98 1723
0 3072 7 1 2 95 1724
0 3073 7 1 2 99 1725
0 3074 7 1 2 96 1726
0 3075 5 10 1 1737
0 3086 5 10 1 1749
0 3097 5 10 1 1763
0 3108 5 10 1 1771
0 3119 5 10 1 1779
0 3130 5 10 1 1787
0 3141 5 1 1 1945
0 3142 5 1 1 1948
0 3143 5 1 1 1951
0 3144 5 1 1 1954
0 3145 5 1 1 1957
0 3146 5 1 1 1960
0 3147 5 10 1 1794
0 3158 5 10 1 1801
0 3169 5 10 1 1808
0 3180 5 10 1 1815
0 3191 9 2 1 1823
0 3194 5 1 1 1933
0 3195 5 1 1 1936
0 3196 5 1 1 1939
0 3197 5 1 1 1942
0 3198 5 1 1 1963
0 3199 5 1 1 1966
0 3200 9 2 1 1474
0 3203 5 1 1 1969
3 3357 9 0 1 2705
3 3358 9 0 1 2706
3 3359 9 0 1 2707
3 3360 9 0 1 2708
0 3401 7 1 3 462 1093 2824
0 3402 7 1 3 473 1094 2826
0 3403 7 1 3 427 1095 2828
0 3404 7 1 3 440 1096 2830
0 3405 7 1 2 1081 2823
0 3406 7 1 2 1082 2825
0 3407 7 1 2 1083 2827
0 3408 7 1 2 1084 2829
0 3409 7 1 3 394 1097 2840
0 3410 7 1 3 405 1098 2842
0 3411 7 1 3 416 1099 2844
0 3412 7 1 3 379 1100 2846
0 3413 7 1 2 1085 2839
0 3414 7 1 2 1086 2841
0 3415 7 1 2 1087 2843
0 3416 7 1 2 1088 2845
0 3444 7 1 2 1281 2902
0 3445 7 1 3 484 1282 2904
0 3446 7 1 3 495 1283 2906
0 3447 7 1 2 1686 2901
0 3448 7 1 2 1687 2903
0 3449 7 1 2 1688 2905
0 3450 7 1 3 508 1101 2914
0 3451 7 1 3 528 1102 2916
0 3452 7 1 3 539 1103 2918
0 3453 7 1 2 1089 2913
0 3454 7 1 2 1090 2915
0 3455 7 1 2 1091 2917
0 3456 7 2 2 2920 2350
0 3459 7 1 3 395 1284 2927
0 3460 7 1 3 406 1285 2929
0 3461 7 1 3 417 1286 2931
0 3462 7 1 3 380 1287 2933
0 3463 7 1 2 1689 2926
0 3464 7 1 2 1690 2928
0 3465 7 1 2 1691 2930
0 3466 7 1 2 1692 2932
0 3481 7 1 3 509 1293 2974
0 3482 5 1 1 2980
0 3483 7 1 3 529 1294 2976
0 3484 7 1 3 540 1295 2978
0 3485 7 1 2 1272 2973
0 3486 7 1 2 1273 2975
0 3487 7 1 2 1274 2977
0 3488 7 1 2 1296 2988
0 3489 7 1 3 485 1297 2990
0 3490 7 1 3 496 1298 2992
0 3491 7 1 2 1275 2987
0 3492 7 1 2 1276 2989
0 3493 7 1 2 1277 2991
0 3502 7 1 2 1299 2999
0 3503 7 1 2 1300 3006
0 3504 7 1 3 463 1288 3016
0 3505 7 1 3 474 1289 3018
0 3506 7 1 3 428 1290 3020
0 3507 7 1 3 441 1291 3022
0 3508 7 1 2 1693 3015
0 3509 7 1 2 1694 3017
0 3510 7 1 2 1695 3019
0 3511 7 1 2 1696 3021
0 3512 6 1 2 1925 3031
0 3513 6 1 2 1922 3032
0 3514 6 1 2 1931 3033
0 3515 6 1 2 1928 3034
0 3558 6 1 2 1949 3141
0 3559 6 1 2 1946 3142
0 3560 6 1 2 1955 3143
0 3561 6 1 2 1952 3144
0 3562 6 1 2 1961 3145
0 3563 6 1 2 1958 3146
3 3604 9 0 1 3192
0 3605 6 1 2 1937 3194
0 3606 6 1 2 1934 3195
0 3607 6 1 2 1943 3196
0 3608 6 1 2 1940 3197
0 3609 6 1 2 1967 3198
0 3610 6 1 2 1964 3199
3 3613 5 0 1 3193
0 3614 7 1 2 2883 2892
0 3615 7 1 2 1484 2893
0 3616 7 1 3 201 2654 1180
0 3617 7 1 3 204 2655 1181
0 3618 7 1 3 198 2656 1182
0 3619 7 1 3 195 2657 1183
0 3620 7 1 3 192 2658 1184
0 3621 7 1 3 183 2682 1204
0 3622 7 1 3 189 2683 1205
0 3623 7 1 3 156 2684 1206
0 3624 7 1 3 150 2685 1207
0 3625 7 1 2 2884 2894
0 3626 7 1 2 1485 2895
0 3627 7 1 3 202 2729 1242
0 3628 7 1 3 205 2730 1243
0 3629 7 1 3 199 2731 1244
0 3630 7 1 3 196 2732 1245
0 3631 7 1 3 193 2733 1246
0 3632 7 1 3 184 2757 1266
0 3633 7 1 3 190 2758 1267
0 3634 7 1 3 157 2759 1268
0 3635 7 1 3 151 2760 1269
0 3636 7 1 2 2885 2896
0 3637 7 1 2 1486 2897
0 3638 7 1 3 110 3076 1750
0 3639 7 1 2 2886 2898
0 3640 7 1 2 1487 2899
0 3641 7 1 3 12 2780 1346
0 3642 7 1 3 111 3042 1716
0 3643 7 1 3 47 3043 1717
0 3644 7 1 3 101 3044 1718
0 3645 7 1 3 92 3045 1719
0 3646 7 1 3 44 3046 1720
0 3647 7 1 3 77 2781 1347
0 3648 7 1 3 74 2782 1348
0 3649 7 1 3 68 2783 1349
0 3650 7 1 3 15 2784 1350
0 3651 7 1 3 48 3077 1751
0 3652 7 1 3 102 3078 1752
0 3653 7 1 3 93 3079 1753
0 3654 7 1 3 45 3080 1754
0 3655 7 1 3 78 2802 1370
0 3656 7 1 3 75 2803 1371
0 3657 7 1 3 69 2804 1372
0 3658 7 1 3 16 2805 1373
0 3659 7 1 3 120 3120 1788
0 3660 7 1 3 13 2806 1374
0 3661 7 1 3 118 3098 1772
0 3662 7 1 3 177 2686 1208
0 3663 7 1 3 178 2761 1270
0 3664 3 1 2 2831 3401
0 3665 3 1 2 2832 3402
0 3666 3 1 2 2833 3403
0 3667 3 1 2 2834 3404
0 3668 3 1 3 2835 3405 464
0 3669 3 1 3 2836 3406 475
0 3670 3 1 3 2837 3407 429
0 3671 3 1 3 2838 3408 442
0 3672 3 1 2 2847 3409
0 3673 3 1 2 2848 3410
0 3674 3 1 2 2849 3411
0 3675 3 1 2 2850 3412
0 3676 3 1 3 2851 3413 396
0 3677 3 1 3 2852 3414 407
0 3678 3 1 3 2853 3415 418
0 3679 3 1 3 2854 3416 381
0 3680 7 1 2 291 2856
0 3681 7 1 2 287 2857
0 3682 7 1 2 279 2858
0 3683 7 1 2 271 2859
0 3684 7 1 2 263 2860
0 3685 7 1 2 240 2862
0 3686 7 1 2 232 2863
0 3687 7 1 2 224 2864
0 3688 7 1 2 216 2865
0 3689 7 1 2 208 2866
0 3691 5 8 1 2900
0 3700 3 1 2 2907 3444
0 3701 3 1 2 2908 3445
0 3702 3 1 2 2909 3446
0 3703 3 1 3 2911 3448 486
0 3704 3 1 3 2912 3449 497
0 3705 3 2 2 2910 3447
0 3708 3 1 2 2919 3450
0 3709 3 1 2 2921 3451
0 3710 3 1 2 2922 3452
0 3711 3 1 3 2923 3453 510
0 3712 3 1 3 2924 3454 530
0 3713 3 1 3 2925 3455 541
0 3715 3 1 2 2934 3459
0 3716 3 1 2 2935 3460
0 3717 3 1 2 2936 3461
0 3718 3 1 2 2937 3462
0 3719 3 1 3 2938 3463 397
0 3720 3 1 3 2939 3464 408
0 3721 3 1 3 2940 3465 419
0 3722 3 1 3 2941 3466 382
0 3723 7 1 2 371 2943
0 3724 7 1 2 365 2944
0 3725 7 1 2 357 2945
0 3726 7 1 2 347 2946
0 3727 7 1 2 330 2949
0 3728 7 1 2 322 2950
0 3729 7 1 2 314 2951
0 3730 7 1 2 306 2952
0 3731 7 1 2 298 2953
0 3732 3 5 2 2947 2958
0 3738 7 1 2 85 2965
0 3739 7 1 2 87 2966
0 3740 7 1 2 35 2967
0 3741 7 1 2 36 2968
0 3742 3 1 2 2979 3481
0 3743 3 1 2 2981 3483
0 3744 3 1 2 2982 3484
0 3745 3 1 3 2983 3485 511
0 3746 3 1 3 2985 3486 531
0 3747 3 1 3 2986 3487 542
0 3748 3 1 2 2993 3488
0 3749 3 1 2 2994 3489
0 3750 3 1 2 2995 3490
0 3751 3 1 3 2997 3492 487
0 3752 3 1 3 2998 3493 498
0 3753 5 1 1 3001
0 3754 5 1 1 3004
0 3755 5 1 1 3008
0 3756 5 1 1 3011
0 3757 3 1 2 3013 3502
0 3758 7 1 3 1325 449 3005
0 3759 3 1 2 3014 3503
0 3760 7 1 3 1326 450 3012
0 3761 7 1 2 1683 3002
0 3762 7 1 2 1684 3009
0 3763 3 1 2 3023 3504
0 3764 3 1 2 3024 3505
0 3765 3 1 2 3025 3506
0 3766 3 1 2 3026 3507
0 3767 3 1 3 3027 3508 465
0 3768 3 1 3 3028 3509 476
0 3769 3 1 3 3029 3510 430
0 3770 3 1 3 3030 3511 443
0 3771 6 3 2 3512 3513
0 3775 6 3 2 3514 3515
0 3779 5 1 1 3036
0 3780 5 1 1 3039
0 3781 7 1 3 117 3099 1773
0 3782 7 1 3 126 3100 1774
0 3783 7 1 3 127 3101 1775
0 3784 7 1 3 128 3102 1776
0 3785 7 1 3 131 3121 1789
0 3786 7 1 3 129 3122 1790
0 3787 7 1 3 119 3123 1791
0 3788 7 1 3 130 3124 1792
0 3789 6 3 2 3558 3559
0 3793 6 3 2 3560 3561
0 3797 6 2 2 3562 3563
0 3800 7 1 3 122 3148 1802
0 3801 7 1 3 113 3149 1803
0 3802 7 1 3 53 3150 1804
0 3803 7 1 3 114 3151 1805
0 3804 7 1 3 115 3152 1806
0 3805 7 1 3 52 3170 1816
0 3806 7 1 3 112 3171 1817
0 3807 7 1 3 116 3172 1818
0 3808 7 1 3 121 3173 1819
0 3809 7 1 3 125 3174 1820
0 3810 6 2 2 3607 3608
0 3813 6 2 2 3605 3606
0 3816 7 2 2 3482 2984
0 3819 3 2 2 2996 3491
0 3822 5 1 1 3201
0 3823 6 1 2 3202 3203
0 3824 6 2 2 3609 3610
0 3827 5 1 1 3457
0 3828 3 1 2 3739 2970
0 3829 3 1 2 3740 2971
0 3830 3 1 2 3741 2972
0 3831 3 1 2 3738 2969
0 3834 5 1 1 3664
0 3835 5 1 1 3665
0 3836 5 1 1 3666
0 3837 5 1 1 3667
0 3838 5 1 1 3672
0 3839 5 1 1 3673
0 3840 5 1 1 3674
0 3841 5 1 1 3675
0 3842 3 6 2 3681 2868
0 3849 3 5 2 3682 2869
0 3855 3 5 2 3683 2870
0 3861 3 5 2 3684 2871
0 3867 3 5 2 3685 2872
0 3873 3 7 2 3686 2873
0 3881 3 5 2 3687 2874
0 3887 3 5 2 3688 2875
0 3893 3 5 2 3689 2876
0 3908 5 1 1 3701
0 3909 5 1 1 3702
0 3911 5 2 1 3700
0 3914 5 1 1 3708
0 3915 5 1 1 3709
0 3916 5 1 1 3710
0 3917 5 1 1 3715
0 3918 5 1 1 3716
0 3919 5 1 1 3717
0 3920 5 1 1 3718
0 3921 3 5 2 3724 2955
0 3927 3 5 2 3725 2956
0 3933 3 5 2 3726 2957
0 3942 3 5 2 3727 2959
0 3948 3 7 2 3728 2960
0 3956 3 5 2 3729 2961
0 3962 3 5 2 3730 2962
0 3968 3 6 2 3731 2963
0 3975 5 1 1 3742
0 3976 5 1 1 3743
0 3977 5 1 1 3744
0 3978 5 1 1 3749
0 3979 5 1 1 3750
0 3980 7 1 3 451 1301 3754
0 3981 7 1 3 452 1302 3756
0 3982 7 1 2 1278 3753
0 3983 7 1 2 1279 3755
0 3984 5 2 1 3757
0 3987 5 1 1 3759
0 3988 5 1 1 3763
0 3989 5 1 1 3764
0 3990 5 1 1 3765
0 3991 5 1 1 3766
0 3998 7 1 3 3458 3125 3131
0 4008 3 2 2 3723 2954
0 4011 3 2 2 3680 2867
0 4021 5 2 1 3748
0 4024 6 1 2 1970 3822
0 4027 5 1 1 3706
0 4031 7 1 2 3828 1584
0 4032 7 1 3 24 2887 3692
0 4033 7 1 3 25 1488 3693
0 4034 7 1 3 26 2888 3694
0 4035 7 1 3 81 1489 3695
0 4036 7 1 2 3829 1585
0 4037 7 1 3 79 2889 3696
0 4038 7 1 3 23 1490 3697
0 4039 7 1 3 82 2890 3698
0 4040 7 1 3 80 1491 3699
0 4041 7 1 2 3830 1586
0 4042 7 1 2 3831 1587
0 4067 7 2 2 3733 521
0 4080 7 3 2 522 3734
0 4088 7 2 2 3834 3668
0 4091 7 2 2 3835 3669
0 4094 7 2 2 3836 3670
0 4097 7 2 2 3837 3671
0 4100 7 2 2 3838 3676
0 4103 7 2 2 3839 3677
0 4106 7 2 2 3840 3678
0 4109 7 2 2 3841 3679
0 4144 7 2 2 3908 3703
0 4147 7 2 2 3909 3704
0 4150 9 2 1 3707
0 4153 7 2 2 3914 3711
0 4156 7 2 2 3915 3712
0 4159 7 2 2 3916 3713
0 4183 3 1 2 3758 3980
0 4184 3 1 2 3760 3981
0 4185 3 1 3 3761 3982 453
0 4186 3 1 3 3762 3983 454
0 4188 5 2 1 3772
0 4191 5 2 1 3776
0 4196 7 1 3 3777 3773 3037
0 4197 7 1 3 3987 3126 3132
0 4198 7 1 2 3920 3722
0 4199 5 1 1 3817
0 4200 5 2 1 3790
0 4203 5 2 1 3794
0 4206 9 2 1 3798
0 4209 9 2 1 3799
0 4212 9 2 1 3735
0 4215 9 2 1 3736
0 4219 9 2 1 3737
0 4223 5 1 1 3811
0 4224 5 1 1 3814
0 4225 7 2 2 3918 3720
0 4228 7 2 2 3919 3721
0 4231 7 2 2 3991 3770
0 4234 7 2 2 3917 3719
0 4237 7 2 2 3989 3768
0 4240 7 2 2 3990 3769
0 4243 7 2 2 3988 3767
0 4246 7 2 2 3976 3746
0 4249 7 2 2 3977 3747
0 4252 7 2 2 3975 3745
0 4255 7 2 2 3978 3751
0 4258 7 2 2 3979 3752
0 4263 5 1 1 3820
0 4264 6 2 2 4024 3823
0 4267 5 1 1 3825
0 4268 7 1 2 455 3894
0 4269 5 1 1 3912
0 4270 5 1 1 3985
0 4271 7 1 2 3895 456
3 4272 5 0 1 4031
0 4273 3 1 4 4032 4033 3614 3615
0 4274 3 1 4 4034 4035 3625 3626
3 4275 5 0 1 4036
0 4276 3 1 4 4037 4038 3636 3637
0 4277 3 1 4 4039 4040 3639 3640
3 4278 5 0 1 4041
3 4279 5 0 1 4042
0 4280 7 3 2 3888 466
0 4284 7 5 2 3882 477
0 4290 7 6 2 431 3874
0 4297 7 1 2 3868 444
0 4298 7 2 2 3862 398
0 4301 7 3 2 3856 409
0 4305 7 4 2 3850 420
0 4310 7 5 2 3843 383
0 4316 7 3 2 467 3889
0 4320 7 4 2 478 3883
0 4325 7 5 2 432 3875
0 4331 7 1 2 445 3869
0 4332 7 3 2 399 3863
0 4336 7 5 2 410 3857
0 4342 7 6 2 421 3851
0 4349 7 7 2 384 3844
0 4357 5 6 1 3969
0 4364 5 10 1 3963
0 4375 9 3 1 3964
0 4379 7 5 2 3957 488
0 4385 7 6 2 499 3949
0 4392 7 1 2 3943 512
0 4396 7 3 2 3934 532
0 4400 7 4 2 3928 543
0 4405 5 6 1 3922
0 4412 9 5 1 3923
0 4418 5 6 1 3970
0 4425 5 10 1 3965
0 4436 9 3 1 3966
0 4440 7 4 2 489 3958
0 4445 7 5 2 500 3950
0 4451 7 1 2 513 3944
0 4456 7 5 2 533 3935
0 4462 7 6 2 544 3929
0 4469 9 7 1 3924
0 4477 5 6 1 3925
0 4512 9 2 1 3971
0 4515 5 1 1 4183
0 4516 5 1 1 4184
0 4521 5 1 1 4009
0 4523 5 1 1 4012
0 4524 5 3 1 4198
0 4532 5 3 1 3986
0 4547 7 1 3 3913 3175 3181
0 4548 9 2 1 3896
0 4551 9 2 1 3890
0 4554 9 2 1 3884
0 4557 9 2 1 3876
0 4560 9 2 1 3870
0 4563 9 2 1 3864
0 4566 9 2 1 3858
0 4569 9 2 1 3852
0 4572 9 2 1 3845
0 4575 4 2 2 433 3877
0 4578 9 2 1 3897
0 4581 9 2 1 3891
0 4584 9 2 1 3885
0 4587 9 2 1 3871
0 4590 9 2 1 3865
0 4593 9 2 1 3859
0 4596 9 2 1 3853
0 4599 9 2 1 3878
0 4602 9 2 1 3846
0 4605 4 2 2 434 3879
0 4608 4 2 2 385 3847
0 4611 9 2 1 3959
0 4614 9 2 1 3951
0 4617 9 2 1 3945
0 4621 9 2 1 3936
0 4624 9 2 1 3930
0 4627 4 2 2 501 3952
0 4630 9 2 1 3960
0 4633 9 2 1 3946
0 4637 9 2 1 3937
0 4640 9 2 1 3931
0 4643 9 2 1 3953
0 4646 4 2 2 502 3954
0 4649 9 2 1 3932
0 4652 9 2 1 3938
0 4655 9 2 1 3926
0 4658 9 2 1 3947
0 4662 9 2 1 3961
0 4665 9 2 1 3955
0 4668 9 2 1 3972
0 4671 9 2 1 3967
0 4674 9 2 1 3880
0 4677 9 2 1 3872
0 4680 9 2 1 3892
0 4683 9 2 1 3886
0 4686 9 2 1 3898
0 4689 9 2 1 3854
0 4692 9 2 1 3848
0 4695 9 2 1 3866
0 4698 9 2 1 3860
0 4701 6 1 2 3815 4223
0 4702 6 1 2 3812 4224
0 4720 5 1 1 4022
0 4721 6 1 2 4023 4263
0 4724 5 1 1 4148
0 4725 5 1 1 4145
0 4726 5 1 1 4160
0 4727 5 1 1 4157
0 4728 5 1 1 4154
0 4729 5 1 1 4098
0 4730 5 1 1 4095
0 4731 5 1 1 4092
0 4732 5 1 1 4089
0 4733 5 1 1 4110
0 4734 5 1 1 4107
0 4735 5 1 1 4104
0 4736 5 1 1 4101
3 4737 7 0 2 4273 2878
3 4738 7 0 2 4274 2879
3 4739 7 0 2 4276 2880
3 4740 7 0 2 4277 2881
0 4741 7 1 3 4151 1760 1756
0 4855 5 1 1 4213
0 4856 6 1 2 4214 2712
0 4908 6 1 2 4216 2718
0 4909 5 1 1 4217
0 4939 7 2 2 4515 4185
0 4942 7 1 2 4516 4186
0 4947 5 1 1 4220
0 4953 7 1 3 4189 3778 3779
0 4954 7 1 3 3774 4192 3780
0 4955 7 1 3 4193 4190 3040
0 4956 7 1 3 4111 3103 3109
0 4957 7 1 3 4108 3104 3110
0 4958 7 1 3 4105 3105 3111
0 4959 7 1 3 4102 3106 3112
0 4960 7 1 3 4161 3127 3133
0 4961 7 1 3 4158 3128 3134
0 4965 5 1 1 4226
0 4966 5 1 1 4229
0 4967 5 1 1 4232
0 4968 5 1 1 4235
0 4972 5 1 1 4247
0 4973 5 1 1 4250
0 4974 5 1 1 4253
0 4975 6 1 2 4254 4199
0 4976 5 1 1 4207
0 4977 5 1 1 4210
0 4978 7 1 3 3795 3791 4208
0 4979 7 1 3 4204 4201 4211
0 4980 7 1 3 4099 3153 3159
0 4981 7 1 3 4096 3154 3160
0 4982 7 1 3 4093 3155 3161
0 4983 7 1 3 4090 3156 3162
0 4984 7 1 3 4155 3176 3182
0 4985 7 1 3 4149 3177 3183
0 4986 7 1 3 4146 3178 3184
0 4987 7 1 3 4152 3179 3185
0 5049 6 2 2 4701 4702
0 5052 5 1 1 4238
0 5053 5 1 1 4241
0 5054 5 1 1 4244
0 5055 5 1 1 4256
0 5056 5 1 1 4259
0 5057 6 1 2 3821 4720
0 5058 5 1 1 4265
0 5059 6 1 2 4266 4267
0 5060 7 1 4 4724 4725 4269 4027
0 5061 7 1 4 4726 4727 3827 4728
0 5062 7 1 4 4729 4730 4731 4732
0 5063 7 1 4 4733 4734 4735 4736
0 5065 7 1 2 4358 4376
0 5066 7 1 3 4365 4359 4380
0 5067 7 1 2 4419 4437
0 5068 7 1 3 4426 4420 4441
0 5069 5 1 1 4549
0 5070 6 1 2 4550 2628
0 5071 5 1 1 4552
0 5072 6 1 2 4553 2629
0 5073 5 1 1 4555
0 5074 6 1 2 4556 2630
0 5075 5 1 1 4558
0 5076 6 1 2 4559 2631
0 5077 5 1 1 4561
0 5078 6 1 2 4562 2632
0 5079 5 1 1 4564
0 5080 6 1 2 4565 2633
0 5081 5 1 1 4567
0 5082 6 1 2 4568 2634
0 5083 5 1 1 4570
0 5084 6 1 2 4571 2635
0 5085 5 1 1 4573
0 5086 6 1 2 4574 2636
0 5087 5 1 1 4576
0 5088 6 1 2 4579 2638
0 5089 5 1 1 4580
0 5090 6 1 2 4582 2639
0 5091 5 1 1 4583
0 5092 6 1 2 4585 2640
0 5093 5 1 1 4586
0 5094 6 1 2 4588 2641
0 5095 5 1 1 4589
0 5096 6 1 2 4591 2642
0 5097 5 1 1 4592
0 5098 6 1 2 4594 2643
0 5099 5 1 1 4595
0 5100 6 1 2 4597 2644
0 5101 5 1 1 4598
0 5102 6 1 2 4600 2645
0 5103 5 1 1 4601
0 5104 6 1 2 4603 2646
0 5105 5 1 1 4604
0 5106 5 1 1 4612
0 5107 6 1 2 4613 2709
0 5108 5 1 1 4615
0 5109 6 1 2 4616 2710
0 5110 5 1 1 4618
0 5111 6 1 2 4619 2711
0 5112 6 1 2 1892 4855
0 5113 5 1 1 4622
0 5114 6 1 2 4623 2713
0 5115 5 1 1 4625
0 5116 6 1 2 4626 2714
0 5117 7 1 2 4366 4381
0 5118 7 1 2 4367 4382
0 5119 7 1 2 56 4406
0 5120 5 1 1 4628
0 5121 6 1 2 4631 2716
0 5122 5 1 1 4632
0 5123 6 1 2 4634 2717
0 5124 5 1 1 4635
0 5125 6 1 2 1910 4909
0 5126 6 1 2 4638 2719
0 5127 5 1 1 4639
0 5128 6 1 2 4641 2720
0 5129 5 1 1 4642
0 5130 6 1 2 4644 2721
0 5131 5 1 1 4645
0 5132 7 1 2 4427 4442
0 5133 7 1 2 4428 4443
0 5135 5 1 1 4650
0 5136 5 1 1 4653
0 5137 6 1 2 4656 4521
0 5138 5 1 1 4657
0 5139 5 1 1 4659
0 5140 6 1 2 4660 4947
0 5141 5 1 1 4675
0 5142 5 1 1 4678
0 5143 5 1 1 4681
0 5144 5 1 1 4684
0 5145 6 1 2 4687 4523
0 5146 5 1 1 4688
0 5147 4 1 2 4953 4196
0 5148 4 1 2 4954 4955
0 5150 5 2 1 4525
0 5153 6 1 2 4230 4965
0 5154 6 1 2 4227 4966
0 5155 6 1 2 4236 4967
0 5156 6 1 2 4233 4968
0 5157 5 2 1 4533
0 5160 6 1 2 4251 4972
0 5161 6 1 2 4248 4973
0 5162 6 1 2 3818 4974
0 5163 7 1 3 4202 3796 4976
0 5164 7 1 3 3792 4205 4977
0 5165 7 1 3 4942 3157 3163
0 5166 5 2 1 4513
0 5169 9 2 1 4291
0 5172 5 1 1 4606
0 5173 9 2 1 4326
0 5176 5 1 1 4609
0 5177 9 2 1 4350
0 5180 9 2 1 4407
0 5183 9 2 1 4360
0 5186 9 2 1 4361
0 5189 9 2 1 4368
0 5192 9 2 1 4369
0 5195 9 2 1 4386
0 5198 5 1 1 4647
0 5199 9 2 1 4421
0 5202 9 2 1 4429
0 5205 9 2 1 4446
0 5208 9 2 1 4422
0 5211 9 2 1 4430
0 5214 9 2 1 4478
0 5217 9 2 1 4470
0 5220 9 2 1 4479
0 5223 5 1 1 4663
0 5224 5 1 1 4666
0 5225 5 1 1 4669
0 5226 5 1 1 4672
0 5227 5 1 1 4690
0 5228 5 1 1 4693
0 5229 5 1 1 4696
0 5230 5 1 1 4699
0 5232 6 1 2 4242 5052
0 5233 6 1 2 4239 5053
0 5234 6 1 2 4260 5055
0 5235 6 1 2 4257 5056
0 5236 6 2 2 4721 5057
0 5239 6 1 2 3826 5058
3 5240 7 0 3 5060 5061 4270
0 5241 5 1 1 4940
0 5242 6 1 2 1826 5069
0 5243 6 1 2 1829 5071
0 5244 6 1 2 1832 5073
0 5245 6 1 2 1835 5075
0 5246 6 1 2 1838 5077
0 5247 6 1 2 1841 5079
0 5248 6 1 2 1844 5081
0 5249 6 1 2 1847 5083
0 5250 6 1 2 1850 5085
0 5252 6 1 2 1856 5089
0 5253 6 1 2 1859 5091
0 5254 6 1 2 1862 5093
0 5255 6 1 2 1865 5095
0 5256 6 1 2 1868 5097
0 5257 6 1 2 1871 5099
0 5258 6 1 2 1874 5101
0 5259 6 1 2 1877 5103
0 5260 6 1 2 1880 5105
0 5261 6 1 2 1883 5106
0 5262 6 1 2 1886 5108
0 5263 6 1 2 1889 5110
0 5264 6 9 2 5112 4856
0 5274 6 1 2 1895 5113
0 5275 6 1 2 1898 5115
0 5282 6 1 2 1904 5122
0 5283 6 1 2 1907 5124
0 5284 6 13 2 4908 5125
0 5298 6 1 2 1913 5127
0 5299 6 1 2 1916 5129
0 5300 6 1 2 1919 5131
0 5303 6 1 2 4654 5135
0 5304 6 1 2 4651 5136
0 5305 6 1 2 4010 5138
0 5306 6 1 2 4221 5139
0 5307 6 1 2 4679 5141
0 5308 6 1 2 4676 5142
0 5309 6 1 2 4685 5143
0 5310 6 1 2 4682 5144
0 5311 6 1 2 4013 5146
0 5312 5 1 1 5050
0 5315 6 3 2 5153 5154
0 5319 6 2 2 5155 5156
0 5324 6 3 2 5160 5161
0 5328 6 2 2 5162 4975
0 5331 4 1 2 5163 4978
0 5332 4 1 2 5164 4979
0 5346 3 2 2 4413 5119
0 5363 6 1 2 4667 5223
0 5364 6 1 2 4664 5224
0 5365 6 1 2 4673 5225
0 5366 6 1 2 4670 5226
0 5367 6 1 2 4694 5227
0 5368 6 1 2 4691 5228
0 5369 6 1 2 4700 5229
0 5370 6 1 2 4697 5230
0 5371 6 2 2 5148 5147
0 5374 9 2 1 4941
0 5377 6 2 2 5232 5233
0 5382 6 2 2 5234 5235
0 5385 6 2 2 5239 5059
3 5388 7 0 3 5062 5063 5241
0 5389 6 6 2 5242 5070
0 5396 6 10 2 5243 5072
0 5407 6 10 2 5244 5074
0 5418 6 5 2 5245 5076
0 5424 6 6 2 5246 5078
0 5431 6 9 2 5247 5080
0 5441 6 10 2 5248 5082
0 5452 6 9 2 5249 5084
0 5462 6 6 2 5250 5086
0 5469 5 1 1 5170
0 5470 6 6 2 5088 5252
0 5477 6 10 2 5090 5253
0 5488 6 9 2 5092 5254
0 5498 6 7 2 5094 5255
0 5506 6 13 2 5096 5256
0 5520 6 15 2 5098 5257
0 5536 6 12 2 5100 5258
0 5549 6 5 2 5102 5259
0 5555 6 6 2 5104 5260
0 5562 6 10 2 5261 5107
0 5573 6 5 2 5262 5109
0 5579 6 6 2 5263 5111
0 5595 6 10 2 5274 5114
0 5606 6 9 2 5275 5116
0 5616 6 1 2 5181 2715
0 5617 5 1 1 5182
0 5618 5 1 1 5184
0 5619 5 1 1 5187
0 5620 5 1 1 5190
0 5621 5 1 1 5193
0 5622 5 1 1 5196
0 5624 6 9 2 5121 5282
0 5634 6 7 2 5123 5283
0 5655 6 15 2 5126 5298
0 5671 6 12 2 5128 5299
0 5684 6 5 2 5130 5300
0 5690 5 1 1 5203
0 5691 5 1 1 5212
0 5692 6 3 2 5303 5304
0 5696 6 3 2 5137 5305
0 5700 6 2 2 5306 5140
0 5703 6 3 2 5307 5308
0 5707 6 3 2 5309 5310
0 5711 6 2 2 5145 5311
0 5726 7 1 2 5167 4514
0 5727 5 1 1 5174
0 5728 5 1 1 5178
0 5730 5 1 1 5200
0 5731 5 1 1 5206
0 5732 5 1 1 5209
0 5733 5 1 1 5215
0 5734 5 1 1 5218
0 5735 5 1 1 5221
0 5736 6 2 2 5365 5366
0 5739 6 2 2 5363 5364
0 5742 6 2 2 5369 5370
0 5745 6 2 2 5367 5368
0 5755 5 1 1 5237
0 5756 6 2 2 5332 5331
0 5954 7 1 2 5265 4397
0 5955 6 1 2 1901 5617
0 5956 5 1 1 5347
0 6005 7 1 2 5285 4457
0 6006 7 1 2 5286 4458
0 6023 5 1 1 5372
0 6024 6 1 2 5373 5312
0 6025 5 2 1 5316
0 6028 5 2 1 5325
0 6031 9 2 1 5320
0 6034 9 2 1 5321
0 6037 9 2 1 5329
0 6040 9 2 1 5330
0 6044 5 1 1 5386
0 6045 3 2 2 5168 5726
0 6048 9 2 1 5266
0 6051 9 2 1 5287
0 6054 9 2 1 5288
0 6065 5 1 1 5375
0 6066 6 1 2 5376 5054
0 6067 5 1 1 5378
0 6068 5 1 1 5383
0 6069 6 1 2 5384 5755
0 6071 7 1 2 5471 4317
0 6072 7 1 3 5478 5472 4321
0 6073 7 1 4 5489 5473 4327 5479
0 6074 7 1 4 5563 4362 4387 4370
0 6075 7 1 2 5390 4281
0 6076 7 1 3 5397 5391 4285
0 6077 7 1 4 5408 5392 4292 5398
0 6078 7 1 4 5625 4423 4447 4431
0 6079 5 1 1 5419
0 6080 7 2 4 5399 5420 5409 5393
0 6083 7 1 2 5400 4286
0 6084 7 1 3 5410 4293 5401
0 6085 7 1 3 5421 5411 5402
0 6086 7 1 2 5403 4287
0 6087 7 1 3 4294 5412 5404
0 6088 7 1 2 5413 4295
0 6089 7 1 2 5422 5414
0 6090 7 1 2 5415 4296
0 6091 7 2 5 5432 5463 5442 5425 5453
0 6094 7 1 2 5426 4299
0 6095 7 1 3 5433 5427 4302
0 6096 7 1 4 5443 5428 4306 5434
0 6097 7 1 5 5454 5444 5429 4311 5435
0 6098 7 1 2 5436 4303
0 6099 7 1 3 5445 4307 5437
0 6100 7 1 4 5455 5446 4312 5438
0 6101 7 1 5 6 5464 5447 5456 5439
0 6102 7 1 2 4308 5448
0 6103 7 1 3 5457 5449 4313
0 6104 7 1 4 7 5465 5450 5458
0 6105 7 1 2 5459 4314
0 6106 7 1 3 8 5466 5460
0 6107 7 1 2 9 5467
0 6108 7 2 4 5550 5490 5480 5474
0 6111 7 1 2 5481 4322
0 6112 7 1 3 5491 4328 5482
0 6113 7 1 3 5551 5492 5483
0 6114 7 1 2 5484 4323
0 6115 7 1 3 5493 4329 5485
0 6116 7 1 2 5494 4330
0 6117 7 2 5 5556 5537 5521 5507 5499
0 6120 7 1 2 5500 4333
0 6121 7 1 3 5508 5501 4337
0 6122 7 1 4 5522 5502 4343 5509
0 6123 7 1 5 5538 5523 5503 4351 5510
0 6124 7 1 2 5511 4338
0 6125 7 1 3 5524 4344 5512
0 6126 7 1 4 5539 5525 4352 5513
0 6127 7 1 4 5557 5526 5514 5540
0 6128 7 1 2 5515 4339
0 6129 7 1 3 5527 4345 5516
0 6130 7 1 4 5541 5528 4353 5517
0 6131 7 1 2 5529 4346
0 6132 7 1 3 5542 5530 4354
0 6133 7 1 3 5558 5531 5543
0 6134 7 1 2 5532 4347
0 6135 7 1 3 5544 5533 4355
0 6136 7 1 2 5545 4356
0 6137 7 1 2 5552 5495
0 6138 7 1 2 5559 5546
0 6139 5 1 1 5574
0 6140 7 2 4 4371 5575 5564 4363
0 6143 7 1 3 5565 4388 4372
0 6144 7 1 3 5576 5566 4373
0 6145 7 1 3 4389 5567 4374
0 6146 7 1 2 5568 4390
0 6147 7 1 2 5577 5569
0 6148 7 1 2 5570 4391
0 6149 7 2 5 5267 4408 5596 5580 5607
0 6152 7 1 2 5581 4068
0 6153 7 1 3 5268 5582 4398
0 6154 7 1 4 5597 5583 4401 5269
0 6155 7 1 5 5608 5598 5584 4414 5270
0 6156 7 1 3 5599 4402 5271
0 6157 7 1 4 5609 5600 4415 5272
0 6158 7 1 5 57 4409 5601 5610 5273
0 6159 7 1 2 4403 5602
0 6160 7 1 3 5611 5603 4416
0 6161 7 1 4 58 4410 5604 5612
0 6162 7 1 2 5613 4417
0 6163 7 1 3 59 4411 5614
0 6164 6 2 2 5616 5955
0 6168 7 2 4 5685 5626 4432 4424
0 6171 7 1 3 5627 4448 4433
0 6172 7 1 3 5686 5628 4434
0 6173 7 1 3 5629 4449 4435
0 6174 7 1 2 5630 4450
0 6175 7 2 5 4480 5672 5656 5289 5635
0 6178 7 1 2 5636 4081
0 6179 7 1 3 5290 5637 4459
0 6180 7 1 4 5657 5638 4463 5291
0 6181 7 1 5 5673 5658 5639 4471 5292
0 6182 7 1 3 5659 4464 5293
0 6183 7 1 4 5674 5660 4472 5294
0 6184 7 1 4 4481 5661 5295 5675
0 6185 7 1 3 5662 4465 5296
0 6186 7 1 4 5676 5663 4473 5297
0 6187 7 1 2 5664 4466
0 6188 7 1 3 5677 5665 4474
0 6189 7 1 3 4482 5666 5678
0 6190 7 1 2 5667 4467
0 6191 7 1 3 5679 5668 4475
0 6192 7 1 2 5680 4476
0 6193 7 1 2 5687 5631
0 6194 7 1 2 4483 5681
0 6197 5 2 1 5693
0 6200 5 2 1 5697
0 6203 5 2 1 5704
0 6206 5 2 1 5708
0 6209 9 2 1 5701
0 6212 9 2 1 5702
0 6215 9 2 1 5712
0 6218 9 2 1 5713
0 6221 6 1 2 5051 6023
0 6234 5 1 1 5757
0 6235 6 1 2 5758 6044
0 6238 9 2 1 5468
0 6241 9 2 1 5394
0 6244 9 2 1 5395
0 6247 9 2 1 5405
0 6250 9 2 1 5406
0 6253 9 2 1 5416
0 6256 9 2 1 5417
0 6259 9 2 1 5430
0 6262 9 2 1 5440
0 6265 9 2 1 5451
0 6268 9 2 1 5461
0 6271 9 2 1 5553
0 6274 9 2 1 5496
0 6277 9 2 1 5475
0 6280 9 2 1 5486
0 6283 9 2 1 5554
0 6286 9 2 1 5497
0 6289 9 2 1 5476
0 6292 9 2 1 5487
0 6295 9 2 1 5560
0 6298 9 2 1 5547
0 6301 9 2 1 5504
0 6304 9 2 1 5534
0 6307 9 2 1 5518
0 6310 9 2 1 5519
0 6313 9 2 1 5561
0 6316 9 2 1 5548
0 6319 9 2 1 5505
0 6322 9 2 1 5535
0 6325 9 2 1 5571
0 6328 9 2 1 5572
0 6331 9 2 1 5585
0 6335 9 2 1 5605
0 6338 9 2 1 5615
0 6341 9 2 1 5688
0 6344 9 2 1 5632
0 6347 9 2 1 5689
0 6350 9 2 1 5633
0 6353 9 2 1 5682
0 6356 9 2 1 5640
0 6359 9 2 1 5669
0 6364 9 2 1 5683
0 6367 9 2 1 5641
0 6370 9 2 1 5670
0 6373 5 1 1 5737
0 6374 5 1 1 5740
0 6375 5 1 1 5743
0 6376 5 1 1 5746
0 6377 6 1 2 4245 6065
0 6378 6 1 2 5238 6068
0 6382 3 1 4 4268 6071 6072 6073
0 6386 3 1 4 3973 5065 5066 6074
0 6388 3 1 4 4271 6075 6076 6077
0 6392 3 1 4 3974 5067 5068 6078
0 6397 3 2 5 4297 6094 6095 6096 6097
0 6411 3 2 2 4324 6116
0 6415 3 3 5 4331 6120 6121 6122 6123
0 6419 3 2 2 4348 6136
0 6427 3 2 5 4392 6152 6153 6154 6155
0 6434 5 1 1 6049
0 6437 3 2 2 4444 6174
0 6441 3 3 5 4451 6178 6179 6180 6181
0 6445 3 2 2 4468 6192
0 6448 5 1 1 6052
0 6449 5 1 1 6055
0 6466 6 2 2 6221 6024
0 6469 5 1 1 6032
0 6470 5 1 1 6035
0 6471 5 1 1 6038
0 6472 5 1 1 6041
0 6473 7 1 3 5317 4526 6033
0 6474 7 1 3 6026 5151 6036
0 6475 7 1 3 5326 4534 6039
0 6476 7 1 3 6029 5158 6042
0 6477 6 1 2 5387 6234
0 6478 6 2 2 6046 133
0 6482 3 2 4 4282 6083 6084 6085
0 6486 4 2 3 4283 6086 6087
0 6490 3 2 3 4288 6088 6089
0 6494 4 2 2 4289 6090
0 6500 3 2 5 4300 6098 6099 6100 6101
0 6504 3 2 4 4304 6102 6103 6104
0 6508 3 2 3 4309 6105 6106
0 6512 3 2 2 4315 6107
0 6516 3 2 4 4318 6111 6112 6113
0 6526 4 2 3 4319 6114 6115
0 6536 3 2 4 4340 6131 6132 6133
0 6539 3 2 5 4334 6124 6125 6126 6127
0 6553 4 2 3 4341 6134 6135
0 6556 4 2 4 4335 6128 6129 6130
0 6566 3 2 4 4377 5117 6143 6144
0 6569 4 2 3 4378 5118 6145
0 6572 3 2 3 4383 6146 6147
0 6575 4 2 2 4384 6148
0 6580 3 2 5 4069 5954 6156 6157 6158
0 6584 3 2 4 4399 6159 6160 6161
0 6587 3 2 3 4404 6162 6163
0 6592 3 2 4 4438 5132 6171 6172
0 6599 4 2 3 4439 5133 6173
0 6606 3 2 4 4460 6187 6188 6189
0 6609 3 2 5 4082 6005 6182 6183 6184
0 6619 4 2 3 4461 6190 6191
0 6622 4 2 4 4083 6006 6185 6186
0 6630 6 1 2 5741 6373
0 6631 6 1 2 5738 6374
0 6632 6 1 2 5747 6375
0 6633 6 1 2 5744 6376
0 6634 6 2 2 6377 6066
0 6637 6 2 2 6069 6378
0 6640 5 1 1 6165
3 6641 7 0 2 6109 6118
3 6643 7 0 2 6141 6150
3 6646 7 0 2 6169 6176
3 6648 7 0 2 6081 6092
0 6650 6 1 2 6239 2637
0 6651 5 1 1 6240
0 6653 5 1 1 6242
0 6655 5 1 1 6245
0 6657 5 1 1 6248
0 6659 5 1 1 6251
0 6660 6 1 2 6254 5087
0 6661 5 1 1 6255
0 6662 6 1 2 6257 5469
0 6663 5 1 1 6258
0 6664 7 1 2 6093 10
0 6666 5 1 1 6260
0 6668 5 1 1 6263
0 6670 5 1 1 6266
0 6672 5 1 1 6269
0 6675 5 1 1 6119
0 6680 5 1 1 6281
0 6681 5 1 1 6293
0 6682 5 1 1 6308
0 6683 5 1 1 6311
0 6689 6 1 2 6326 5120
0 6690 5 1 1 6327
0 6691 6 1 2 6329 5622
0 6692 5 1 1 6330
0 6693 7 1 2 6151 60
0 6695 5 1 1 6332
0 6698 5 1 1 6336
0 6699 6 1 2 6339 5956
0 6700 5 1 1 6340
0 6703 5 1 1 6177
0 6708 5 1 1 6210
0 6709 5 1 1 6213
0 6710 5 1 1 6216
0 6711 5 1 1 6219
0 6712 7 1 3 5698 5694 6211
0 6713 7 1 3 6201 6198 6214
0 6714 7 1 3 5709 5705 6217
0 6715 7 1 3 6207 6204 6220
3 6716 9 0 1 6467
0 6718 7 1 3 6166 1780 3135
0 6719 7 1 3 5152 5318 6469
0 6720 7 1 3 4527 6027 6470
0 6721 7 1 3 5159 5327 6471
0 6722 7 1 3 4535 6030 6472
0 6724 6 2 2 6477 6235
0 6739 5 1 1 6272
0 6740 5 1 1 6275
0 6741 5 1 1 6278
0 6744 5 1 1 6284
0 6745 5 1 1 6287
0 6746 5 1 1 6290
0 6751 5 1 1 6296
0 6752 5 1 1 6299
0 6753 5 1 1 6302
0 6754 5 1 1 6305
0 6755 5 1 1 6323
0 6760 5 1 1 6314
0 6761 5 1 1 6317
0 6762 5 1 1 6320
0 6772 5 1 1 6342
0 6773 5 1 1 6345
0 6776 5 1 1 6348
0 6777 5 1 1 6351
0 6782 5 1 1 6354
0 6783 5 1 1 6357
0 6784 5 1 1 6360
0 6785 5 1 1 6371
0 6790 5 1 1 6365
0 6791 5 1 1 6368
0 6792 6 2 2 6630 6631
0 6795 6 2 2 6632 6633
0 6801 7 1 2 6110 6416
0 6802 7 1 2 6428 6142
0 6803 7 1 2 6398 6082
0 6804 7 1 2 6170 6442
0 6805 5 1 1 6468
0 6806 6 1 2 1853 6651
0 6807 5 1 1 6483
0 6808 6 1 2 6484 6653
0 6809 5 1 1 6487
0 6810 6 1 2 6488 6655
0 6811 5 1 1 6491
0 6812 6 1 2 6492 6657
0 6813 5 1 1 6495
0 6814 6 1 2 6496 6659
0 6815 6 1 2 4577 6661
0 6816 6 1 2 5171 6663
0 6817 3 5 2 6399 6664
0 6823 5 1 1 6501
0 6824 6 1 2 6502 6666
0 6825 5 1 1 6505
0 6826 6 1 2 6506 6668
0 6827 5 1 1 6509
0 6828 6 1 2 6510 6670
0 6829 5 1 1 6513
0 6830 6 1 2 6514 6672
0 6831 5 2 1 6417
0 6834 5 1 1 6567
0 6835 6 1 2 6568 5618
0 6836 5 1 1 6570
0 6837 6 1 2 6571 5619
0 6838 5 1 1 6573
0 6839 6 1 2 6574 5620
0 6840 5 1 1 6576
0 6841 6 1 2 6577 5621
0 6842 6 1 2 4629 6690
0 6843 6 1 2 5197 6692
0 6844 3 5 2 6429 6693
0 6850 5 1 1 6581
0 6851 6 1 2 6582 6695
0 6852 5 1 1 6585
0 6853 6 1 2 6586 6434
0 6854 5 1 1 6588
0 6855 6 1 2 6589 6698
0 6856 6 1 2 5348 6700
0 6857 5 2 1 6443
0 6860 7 1 3 6199 5699 6708
0 6861 7 1 3 5695 6202 6709
0 6862 7 1 3 6205 5710 6710
0 6863 7 1 3 5706 6208 6711
0 6866 3 5 3 4197 6718 3785
0 6872 4 1 2 6719 6473
0 6873 4 1 2 6720 6474
0 6874 4 1 2 6721 6475
0 6875 4 1 2 6722 6476
0 6876 5 1 1 6638
3 6877 9 0 1 6725
0 6879 7 1 2 6047 6479
0 6880 7 1 2 6480 134
0 6881 3 2 2 6412 6137
0 6884 5 1 1 6517
0 6885 5 2 1 6413
0 6888 5 1 1 6527
0 6889 5 1 1 6537
0 6890 6 1 2 6538 5176
0 6891 3 2 2 6420 6138
0 6894 5 1 1 6540
0 6895 5 1 1 6554
0 6896 6 1 2 6555 5728
0 6897 5 2 1 6421
0 6900 5 1 1 6557
0 6901 3 2 2 6438 6193
0 6904 5 1 1 6593
0 6905 5 2 1 6439
0 6908 5 1 1 6600
0 6909 3 2 2 6446 6194
0 6912 5 1 1 6607
0 6913 5 1 1 6610
0 6914 5 1 1 6620
0 6915 6 1 2 6621 5734
0 6916 5 2 1 6447
0 6919 5 1 1 6623
0 6922 5 1 1 6635
0 6923 6 1 2 6636 6067
3 6924 3 0 2 6382 6801
3 6925 3 0 2 6386 6802
3 6926 3 0 2 6388 6803
3 6927 3 0 2 6392 6804
0 6930 5 1 1 6726
0 6932 6 2 2 6650 6806
0 6935 6 1 2 6243 6807
0 6936 6 1 2 6246 6809
0 6937 6 1 2 6249 6811
0 6938 6 1 2 6252 6813
0 6939 6 1 2 6660 6815
0 6940 6 1 2 6662 6816
0 6946 6 1 2 6261 6823
0 6947 6 1 2 6264 6825
0 6948 6 1 2 6267 6827
0 6949 6 1 2 6270 6829
0 6953 6 1 2 5185 6834
0 6954 6 1 2 5188 6836
0 6955 6 1 2 5191 6838
0 6956 6 1 2 5194 6840
0 6957 6 1 2 6689 6842
0 6958 6 1 2 6691 6843
0 6964 6 1 2 6333 6850
0 6965 6 1 2 6050 6852
0 6966 6 1 2 6337 6854
0 6967 6 2 2 6699 6856
0 6973 4 1 2 6860 6712
0 6974 4 1 2 6861 6713
0 6975 4 1 2 6862 6714
0 6976 4 1 2 6863 6715
0 6977 5 1 1 6793
0 6978 5 1 1 6796
0 6979 3 3 2 6879 6880
0 6987 6 1 2 4610 6889
0 6990 6 1 2 5179 6895
0 6999 6 1 2 5219 6914
0 7002 6 1 2 5379 6922
0 7003 6 2 2 6873 6872
0 7006 6 2 2 6875 6874
0 7011 7 1 3 6867 2687 2693
0 7012 7 1 3 6868 2762 2768
0 7013 7 1 3 6869 2785 2791
3 7015 5 0 1 6870
0 7016 7 1 3 6871 2807 2813
0 7018 6 1 2 6935 6808
0 7019 6 1 2 6936 6810
0 7020 6 1 2 6937 6812
0 7021 6 1 2 6938 6814
0 7022 5 1 1 6939
0 7023 5 4 1 6818
0 7028 6 2 2 6946 6824
0 7031 6 2 2 6947 6826
0 7034 6 2 2 6948 6828
0 7037 6 2 2 6949 6830
0 7040 7 1 2 6819 6079
0 7041 7 2 2 6832 6675
0 7044 6 1 2 6953 6835
0 7045 6 1 2 6954 6837
0 7046 6 1 2 6955 6839
0 7047 6 1 2 6956 6841
0 7048 5 1 1 6957
0 7049 5 4 1 6845
0 7054 6 2 2 6964 6851
0 7057 6 2 2 6965 6853
0 7060 6 2 2 6966 6855
0 7064 7 1 2 6846 6139
0 7065 7 2 2 6858 6703
0 7072 5 1 1 6882
0 7073 6 1 2 6883 5172
0 7074 5 1 1 6886
0 7075 6 1 2 6887 5727
0 7076 6 2 2 6890 6987
0 7079 5 1 1 6892
0 7080 6 2 2 6896 6990
0 7083 5 1 1 6898
0 7084 5 1 1 6902
0 7085 6 1 2 6903 5198
0 7086 5 1 1 6906
0 7087 6 1 2 6907 5731
0 7088 5 1 1 6910
0 7089 6 1 2 6911 6912
0 7090 6 2 2 6915 6999
0 7093 5 1 1 6917
0 7094 6 2 2 6974 6973
0 7097 6 2 2 6976 6975
0 7101 6 2 2 7002 6923
0 7105 5 1 1 6933
0 7110 5 1 1 6968
0 7114 7 1 3 6980 605 1757
0 7115 5 1 1 7019
0 7116 5 1 1 7021
0 7125 7 1 2 6820 7018
0 7126 7 1 2 6821 7020
0 7127 7 1 2 6822 7022
0 7130 5 1 1 7045
0 7131 5 1 1 7047
0 7139 7 1 2 6847 7044
0 7140 7 1 2 6848 7046
0 7141 7 1 2 6849 7048
0 7146 7 1 3 6934 1764 3113
0 7147 7 1 3 6969 1781 3136
0 7149 5 1 1 7004
0 7150 5 1 1 7007
0 7151 6 1 2 7008 6876
0 7152 6 1 2 4607 7072
0 7153 6 1 2 5175 7074
0 7158 6 1 2 4648 7084
0 7159 6 1 2 5207 7086
0 7160 6 1 2 6608 7088
0 7166 5 1 1 7038
0 7167 5 1 1 7035
0 7168 5 1 1 7032
0 7169 5 1 1 7029
0 7170 5 1 1 7061
0 7171 5 1 1 7058
0 7172 5 1 1 7055
0 7173 7 1 2 7115 7024
0 7174 7 1 2 7116 7025
0 7175 7 1 2 6940 7026
0 7176 7 1 2 5423 7027
0 7177 5 1 1 7042
0 7178 7 1 2 7130 7050
0 7179 7 1 2 7131 7051
0 7180 7 1 2 6958 7052
0 7181 7 1 2 5578 7053
0 7182 5 1 1 7066
0 7183 5 1 1 7095
0 7184 6 1 2 7096 6977
0 7185 5 1 1 7098
0 7186 6 1 2 7099 6978
0 7187 7 1 3 7039 1765 3114
0 7188 7 1 3 7036 1766 3115
0 7189 7 1 3 7033 1767 3116
0 7190 3 5 3 4956 7146 3781
0 7196 7 1 3 7062 1782 3137
0 7197 7 1 3 7059 1783 3138
0 7198 3 5 3 4960 7147 3786
0 7204 6 1 2 7102 7149
0 7205 5 1 1 7103
0 7206 6 1 2 6639 7150
0 7207 7 1 3 7030 1795 3164
0 7208 7 1 3 7056 1809 3186
0 7209 6 2 2 7073 7152
0 7212 6 2 2 7075 7153
0 7215 5 1 1 7077
0 7216 6 1 2 7078 7079
0 7217 5 1 1 7081
0 7218 6 1 2 7082 7083
0 7219 6 2 2 7085 7158
0 7222 6 2 2 7087 7159
0 7225 6 2 2 7089 7160
0 7228 5 1 1 7091
0 7229 6 1 2 7092 7093
0 7236 3 2 2 7173 7125
0 7239 3 2 2 7174 7126
0 7242 3 2 2 7175 7127
0 7245 3 2 2 7176 7040
0 7250 3 6 2 7178 7139
0 7257 3 2 2 7179 7140
0 7260 3 2 2 7180 7141
0 7263 3 2 2 7181 7064
0 7268 6 1 2 6794 7183
0 7269 6 1 2 6797 7185
0 7270 3 5 3 4957 7187 3782
0 7276 3 5 3 4958 7188 3783
0 7282 3 5 3 4959 7189 3784
0 7288 3 5 3 4961 7196 3787
0 7294 3 5 3 3998 7197 3788
0 7300 6 1 2 7005 7205
0 7301 6 2 2 7206 7151
0 7304 3 5 3 4980 7207 3800
0 7310 3 5 3 4984 7208 3805
0 7320 6 1 2 6893 7215
0 7321 6 1 2 6899 7217
0 7328 6 1 2 6918 7228
0 7338 7 1 3 7191 1192 2694
0 7339 7 1 3 7199 2688 2695
0 7340 7 1 3 7192 1254 2769
0 7341 7 1 3 7200 2763 2770
0 7342 7 1 3 7193 1334 2792
0 7349 7 1 3 7201 2786 2793
0 7357 7 1 3 7202 2808 2814
3 7363 5 0 1 7203
0 7364 7 1 3 7194 1358 2815
3 7365 5 0 1 7195
0 7394 6 2 2 7268 7184
0 7397 6 2 2 7269 7186
0 7402 6 2 2 7204 7300
0 7405 5 1 1 7210
0 7406 6 1 2 7211 6884
0 7407 5 1 1 7213
0 7408 6 1 2 7214 6888
0 7409 6 2 2 7320 7216
0 7412 6 2 2 7321 7218
0 7415 5 1 1 7220
0 7416 6 1 2 7221 6904
0 7417 5 1 1 7223
0 7418 6 1 2 7224 6908
0 7419 5 1 1 7226
0 7420 6 1 2 7227 6913
0 7421 6 2 2 7328 7229
0 7424 5 1 1 7246
0 7425 5 1 1 7243
0 7426 5 1 1 7240
0 7427 5 1 1 7237
0 7428 5 1 1 7264
0 7429 5 1 1 7261
0 7430 5 1 1 7258
0 7431 5 1 1 7251
3 7432 5 0 1 7252
0 7433 7 1 3 7311 2659 2665
0 7434 7 1 3 7305 1168 2666
0 7435 3 1 4 7011 7338 3621 2591
0 7436 7 1 3 7271 1193 2696
0 7437 7 1 3 7289 2689 2697
0 7438 7 1 3 7277 1194 2698
0 7439 7 1 3 7295 2690 2699
0 7440 7 1 3 7283 1195 2700
0 7441 7 1 3 7312 2734 2740
0 7442 7 1 3 7306 1230 2741
0 7443 3 1 4 7012 7340 3632 2600
0 7444 7 1 3 7272 1255 2771
0 7445 7 1 3 7290 2764 2772
0 7446 7 1 3 7278 1256 2773
0 7447 7 1 3 7296 2765 2774
0 7448 7 1 3 7284 1257 2775
3 7449 3 0 4 7013 7342 3641 2605
0 7450 7 1 3 7313 3047 3053
0 7451 7 1 3 7307 1704 3054
0 7452 7 1 3 7297 2787 2794
0 7453 7 1 3 7285 1335 2795
0 7454 7 1 3 7291 2788 2796
0 7455 7 1 3 7279 1336 2797
0 7456 7 1 3 7273 1337 2798
0 7457 7 1 3 7314 3081 3087
0 7458 7 1 3 7308 1738 3088
0 7459 7 1 3 7298 2809 2816
0 7460 7 1 3 7286 1359 2817
0 7461 7 1 3 7292 2810 2818
0 7462 7 1 3 7280 1360 2819
0 7463 7 1 3 7274 1361 2820
0 7464 7 1 3 7253 606 602
3 7465 5 0 1 7315
3 7466 5 0 1 7299
3 7467 5 0 1 7293
0 7468 5 1 1 7302
3 7469 3 0 4 7016 7364 3660 2626
3 7470 5 0 1 7309
3 7471 5 0 1 7287
3 7472 5 0 1 7281
3 7473 5 0 1 7275
3 7474 9 0 1 7395
3 7476 9 0 1 7398
0 7479 7 1 2 7303 3069
0 7481 7 1 3 7247 1796 3165
0 7482 7 1 3 7244 1797 3166
0 7483 7 1 3 7241 1798 3167
0 7484 7 1 3 7238 1799 3168
0 7485 7 1 3 7265 1810 3187
0 7486 7 1 3 7262 1811 3188
0 7487 7 1 3 7259 1812 3189
0 7488 7 1 3 7254 1813 3190
0 7489 6 2 2 6981 7255
0 7492 6 1 2 6518 7405
0 7493 6 1 2 6528 7407
0 7498 6 1 2 6594 7415
0 7499 6 1 2 6601 7417
0 7500 6 1 2 6611 7419
3 7503 7 0 9 7105 7166 7167 7168 7169 7424 7425 7426 7427
3 7504 7 0 9 6640 7110 7170 7171 7172 7428 7429 7430 7431
0 7505 3 1 4 7433 7434 3616 2585
3 7506 7 0 2 7435 2676
0 7507 3 1 4 7339 7436 3622 2592
0 7508 3 1 4 7437 7438 3623 2593
0 7509 3 1 4 7439 7440 3624 2594
0 7510 3 1 4 7441 7442 3627 2595
3 7511 7 0 2 7443 2751
0 7512 3 1 4 7341 7444 3633 2601
0 7513 3 1 4 7445 7446 3634 2602
0 7514 3 1 4 7447 7448 3635 2603
3 7515 3 0 4 7450 7451 3646 2610
3 7516 3 0 4 7452 7453 3647 2611
3 7517 3 0 4 7454 7455 3648 2612
3 7518 3 0 4 7349 7456 3649 2613
3 7519 3 0 4 7457 7458 3654 2618
3 7520 3 0 4 7459 7460 3655 2619
3 7521 3 0 4 7461 7462 3656 2620
3 7522 3 0 4 7357 7463 3657 2621
0 7525 3 1 4 4741 7114 2624 7464
0 7526 7 1 3 7468 3129 3139
0 7527 5 1 1 7396
0 7528 5 1 1 7399
0 7529 5 1 1 7403
0 7530 7 1 2 7404 3070
0 7531 3 5 3 4981 7481 3801
0 7537 3 5 3 4982 7482 3802
0 7543 3 5 3 4983 7483 3803
0 7549 3 5 3 5165 7484 3804
0 7555 3 5 3 4985 7485 3806
0 7561 3 5 3 4986 7486 3807
0 7567 3 5 3 4547 7487 3808
0 7573 3 5 3 4987 7488 3809
0 7579 6 2 2 7492 7406
0 7582 6 2 2 7493 7408
0 7585 5 1 1 7410
0 7586 6 1 2 7411 6894
0 7587 5 1 1 7413
0 7588 6 1 2 7414 6900
0 7589 6 2 2 7498 7416
0 7592 6 2 2 7499 7418
0 7595 6 2 2 7500 7420
0 7598 5 1 1 7422
0 7599 6 1 2 7423 6919
3 7600 7 0 2 7505 2648
3 7601 7 0 2 7507 2677
3 7602 7 0 2 7508 2678
3 7603 7 0 2 7509 2679
3 7604 7 0 2 7510 2723
3 7605 7 0 2 7512 2752
3 7606 7 0 2 7513 2753
3 7607 7 0 2 7514 2754
0 7624 7 1 2 6982 7490
0 7625 7 1 2 7491 7256
3 7626 7 0 2 1149 7525
0 7631 7 1 5 565 7527 7528 6805 6930
0 7636 7 1 3 7529 3107 3117
0 7657 6 1 2 6541 7585
0 7658 6 1 2 6558 7587
0 7665 6 1 2 6624 7598
0 7666 7 1 3 7556 2660 2667
0 7667 7 1 3 7532 1169 2668
0 7668 7 1 3 7562 2661 2669
0 7669 7 1 3 7538 1170 2670
0 7670 7 1 3 7568 2662 2671
0 7671 7 1 3 7544 1171 2672
0 7672 7 1 3 7574 2663 2673
0 7673 7 1 3 7550 1172 2674
0 7674 7 1 3 7557 2735 2742
0 7675 7 1 3 7533 1231 2743
0 7676 7 1 3 7563 2736 2744
0 7677 7 1 3 7539 1232 2745
0 7678 7 1 3 7569 2737 2746
0 7679 7 1 3 7545 1233 2747
0 7680 7 1 3 7575 2738 2748
0 7681 7 1 3 7551 1234 2749
0 7682 7 1 3 7576 3082 3089
0 7683 7 1 3 7552 1739 3090
0 7684 7 1 3 7577 3048 3055
0 7685 7 1 3 7553 1705 3056
0 7686 7 1 3 7570 3049 3057
0 7687 7 1 3 7546 1706 3058
0 7688 7 1 3 7564 3050 3059
0 7689 7 1 3 7540 1707 3060
0 7690 7 1 3 7558 3051 3061
0 7691 7 1 3 7534 1708 3062
0 7692 7 1 3 7571 3083 3091
0 7693 7 1 3 7547 1740 3092
0 7694 7 1 3 7565 3084 3093
0 7695 7 1 3 7541 1741 3094
0 7696 7 1 3 7559 3085 3095
0 7697 7 1 3 7535 1742 3096
3 7698 3 0 2 7624 7625
3 7699 5 0 1 7578
3 7700 5 0 1 7572
3 7701 5 0 1 7566
3 7702 5 0 1 7560
3 7703 7 0 3 1156 7631 247
3 7704 5 0 1 7554
3 7705 5 0 1 7548
3 7706 5 0 1 7542
3 7707 5 0 1 7536
0 7708 5 1 1 7580
0 7709 6 1 2 7581 6739
0 7710 5 1 1 7583
0 7711 6 1 2 7584 6744
0 7712 6 2 2 7657 7586
0 7715 6 2 2 7658 7588
0 7718 5 1 1 7590
0 7719 6 1 2 7591 6772
0 7720 5 1 1 7593
0 7721 6 1 2 7594 6776
0 7722 5 1 1 7596
0 7723 6 1 2 7597 5733
0 7724 6 2 2 7665 7599
0 7727 3 1 4 7666 7667 3617 2586
0 7728 3 1 4 7668 7669 3618 2587
0 7729 3 1 4 7670 7671 3619 2588
0 7730 3 1 4 7672 7673 3620 2589
0 7731 3 1 4 7674 7675 3628 2596
0 7732 3 1 4 7676 7677 3629 2597
0 7733 3 1 4 7678 7679 3630 2598
0 7734 3 1 4 7680 7681 3631 2599
3 7735 3 0 4 7682 7683 3638 2604
3 7736 3 0 4 7684 7685 3642 2606
3 7737 3 0 4 7686 7687 3643 2607
3 7738 3 0 4 7688 7689 3644 2608
3 7739 3 0 4 7690 7691 3645 2609
3 7740 3 0 4 7692 7693 3651 2615
3 7741 3 0 4 7694 7695 3652 2616
3 7742 3 0 4 7696 7697 3653 2617
0 7743 6 1 2 6273 7708
0 7744 6 1 2 6285 7710
0 7749 6 1 2 6343 7718
0 7750 6 1 2 6349 7720
0 7751 6 1 2 5216 7722
3 7754 7 0 2 7727 2649
3 7755 7 0 2 7728 2650
3 7756 7 0 2 7729 2651
3 7757 7 0 2 7730 2652
3 7758 7 0 2 7731 2724
3 7759 7 0 2 7732 2725
3 7760 7 0 2 7733 2726
3 7761 7 0 2 7734 2727
0 7762 6 2 2 7743 7709
0 7765 6 2 2 7744 7711
0 7768 5 1 1 7713
0 7769 6 1 2 7714 6751
0 7770 5 1 1 7716
0 7771 6 1 2 7717 6760
0 7772 6 2 2 7749 7719
0 7775 6 2 2 7750 7721
0 7778 6 2 2 7751 7723
0 7781 5 1 1 7725
0 7782 6 1 2 7726 5735
0 7787 6 1 2 6297 7768
0 7788 6 1 2 6315 7770
0 7795 6 1 2 5222 7781
0 7796 5 1 1 7763
0 7797 6 1 2 7764 6740
0 7798 5 1 1 7766
0 7799 6 1 2 7767 6745
0 7800 6 2 2 7787 7769
0 7803 6 2 2 7788 7771
0 7806 5 1 1 7773
0 7807 6 1 2 7774 6773
0 7808 5 1 1 7776
0 7809 6 1 2 7777 6777
0 7810 5 1 1 7779
0 7811 6 1 2 7780 6782
0 7812 6 2 2 7795 7782
0 7815 6 1 2 6276 7796
0 7816 6 1 2 6288 7798
0 7821 6 1 2 6346 7806
0 7822 6 1 2 6352 7808
0 7823 6 1 2 6355 7810
0 7826 6 2 2 7815 7797
0 7829 6 2 2 7816 7799
0 7832 5 1 1 7801
0 7833 6 1 2 7802 6752
0 7834 5 1 1 7804
0 7835 6 1 2 7805 6761
0 7836 6 2 2 7821 7807
0 7839 6 2 2 7822 7809
0 7842 6 2 2 7823 7811
0 7845 5 1 1 7813
0 7846 6 1 2 7814 6790
0 7851 6 1 2 6300 7832
0 7852 6 1 2 6318 7834
0 7859 6 1 2 6366 7845
0 7860 5 1 1 7827
0 7861 6 1 2 7828 6741
0 7862 5 1 1 7830
0 7863 6 1 2 7831 6746
0 7864 6 2 2 7851 7833
0 7867 6 2 2 7852 7835
0 7870 5 1 1 7837
0 7871 6 1 2 7838 5730
0 7872 5 1 1 7840
0 7873 6 1 2 7841 5732
0 7874 5 1 1 7843
0 7875 6 1 2 7844 6783
0 7876 6 2 2 7859 7846
0 7879 6 1 2 6279 7860
0 7880 6 1 2 6291 7862
0 7885 6 1 2 5201 7870
0 7886 6 1 2 5210 7872
0 7887 6 1 2 6358 7874
0 7890 6 2 2 7879 7861
0 7893 6 2 2 7880 7863
0 7896 5 1 1 7865
0 7897 6 1 2 7866 6753
0 7898 5 1 1 7868
0 7899 6 1 2 7869 6762
0 7900 6 2 2 7885 7871
0 7903 6 2 2 7886 7873
0 7906 6 2 2 7887 7875
0 7909 5 1 1 7877
0 7910 6 1 2 7878 6791
0 7917 6 1 2 6303 7896
0 7918 6 1 2 6321 7898
0 7923 6 1 2 6369 7909
0 7924 5 1 1 7891
0 7925 6 1 2 7892 6680
0 7926 5 1 1 7894
0 7927 6 1 2 7895 6681
0 7928 5 1 1 7901
0 7929 6 1 2 7902 5690
0 7930 5 1 1 7904
0 7931 6 1 2 7905 5691
0 7932 6 2 2 7917 7897
0 7935 6 2 2 7918 7899
0 7938 5 1 1 7907
0 7939 6 1 2 7908 6784
0 7940 6 2 2 7923 7910
0 7943 6 1 2 6282 7924
0 7944 6 1 2 6294 7926
0 7945 6 1 2 5204 7928
0 7946 6 1 2 5213 7930
0 7951 6 1 2 6361 7938
0 7954 6 2 2 7943 7925
0 7957 6 2 2 7944 7927
0 7960 6 2 2 7945 7929
0 7963 6 2 2 7946 7931
0 7966 5 1 1 7933
0 7967 6 1 2 7934 6754
0 7968 5 1 1 7936
0 7969 6 1 2 7937 6755
0 7970 6 2 2 7951 7939
0 7973 5 1 1 7941
0 7974 6 1 2 7942 6785
0 7984 6 1 2 6306 7966
0 7985 6 1 2 6324 7968
0 7987 6 1 2 6372 7973
0 7988 7 1 3 7958 6833 1158
0 7989 7 1 3 7955 6418 1159
0 7990 7 1 3 7959 7043 568
0 7991 7 1 3 7956 7177 569
0 7992 5 1 1 7971
0 7993 6 1 2 7972 6448
0 7994 7 1 3 7964 6859 1220
0 7995 7 1 3 7961 6444 1221
0 7996 7 1 3 7965 7067 585
0 7997 7 1 3 7962 7182 586
0 7998 6 2 2 7984 7967
0 8001 6 2 2 7985 7969
0 8004 6 2 2 7987 7974
0 8009 6 1 2 6053 7992
0 8013 3 2 4 7988 7989 7990 7991
0 8017 3 2 4 7994 7995 7996 7997
0 8020 5 1 1 7999
0 8021 6 1 2 8000 6682
0 8022 5 1 1 8002
0 8023 6 1 2 8003 6683
0 8025 6 1 2 8009 7993
0 8026 5 1 1 8005
0 8027 6 1 2 8006 6449
0 8031 6 1 2 6309 8020
0 8032 6 1 2 6312 8022
0 8033 5 1 1 8014
0 8034 6 1 2 6056 8026
0 8035 7 1 2 587 8025
0 8036 5 1 1 8018
0 8037 6 1 2 8031 8021
0 8038 6 1 2 8032 8023
0 8039 6 1 2 8034 8027
0 8040 5 1 1 8038
0 8041 7 1 2 570 8037
0 8042 5 1 1 8039
0 8043 7 1 2 8040 1160
0 8044 7 1 2 8042 1222
0 8045 3 2 2 8043 8041
0 8048 3 2 2 8044 8035
0 8055 6 1 2 8046 8033
0 8056 5 1 1 8047
0 8057 6 1 2 8049 8036
0 8058 5 1 1 8050
0 8059 6 1 2 8015 8056
0 8060 6 1 2 8019 8058
0 8061 6 2 2 8055 8059
0 8064 6 2 2 8057 8060
0 8071 7 1 3 8065 1784 3140
0 8072 7 1 3 8062 1768 3118
0 8073 5 1 1 8063
0 8074 5 1 1 8066
3 8075 3 0 4 7526 8071 3659 2625
3 8076 3 0 4 7636 8072 3661 2627
0 8077 7 1 2 8073 1729
0 8078 7 1 2 8074 1730
0 8079 3 2 2 7530 8077
0 8082 3 2 2 7479 8078
0 8089 7 1 2 8080 3064
0 8090 7 1 2 8083 3065
0 8091 7 1 2 8081 3066
0 8092 7 1 2 8084 3067
0 8093 3 2 2 8089 3071
0 8096 3 2 2 8090 3072
0 8099 3 2 2 8091 3073
0 8102 3 2 2 8092 3074
0 8113 7 1 3 8103 2789 2799
0 8114 7 1 3 8100 1338 2800
0 8115 7 1 3 8104 2811 2821
0 8116 7 1 3 8101 1362 2822
0 8117 7 1 3 8097 2691 2701
0 8118 7 1 3 8094 1196 2702
0 8119 7 1 3 8098 2766 2776
0 8120 7 1 3 8095 1258 2777
0 8121 3 1 4 8117 8118 3662 2703
0 8122 3 1 4 8119 8120 3663 2778
3 8123 3 0 4 8113 8114 3650 2614
3 8124 3 0 4 8115 8116 3658 2622
0 8125 7 1 2 8121 2680
0 8126 7 1 2 8122 2755
3 8127 5 0 1 8125
3 8128 5 0 1 8126
2 2 1 1
2 3 1 1
2 5 1 4
2 6 1 4
2 7 1 4
2 8 1 4
2 9 1 4
2 10 1 4
2 12 1 11
2 13 1 11
2 15 1 14
2 16 1 14
2 18 1 17
2 19 1 17
2 21 1 20
2 22 1 20
2 28 1 27
2 29 1 27
2 30 1 27
2 32 1 31
2 33 1 31
2 35 1 34
2 36 1 34
2 38 1 37
2 39 1 37
2 41 1 40
2 42 1 40
2 44 1 43
2 45 1 43
2 47 1 46
2 48 1 46
2 50 1 49
2 51 1 49
2 55 1 54
2 56 1 54
2 57 1 54
2 58 1 54
2 59 1 54
2 60 1 54
2 62 1 61
2 63 1 61
2 65 1 64
2 66 1 64
2 68 1 67
2 69 1 67
2 71 1 70
2 72 1 70
2 74 1 73
2 75 1 73
2 77 1 76
2 78 1 76
2 84 1 83
2 85 1 83
2 89 1 88
2 90 1 88
2 92 1 91
2 93 1 91
2 95 1 94
2 96 1 94
2 98 1 97
2 99 1 97
2 101 1 100
2 102 1 100
2 104 1 103
2 105 1 103
2 107 1 106
2 108 1 106
2 110 1 109
2 111 1 109
2 124 1 123
2 125 1 123
2 133 1 132
2 134 1 132
2 138 1 137
2 139 1 137
2 142 1 141
2 143 1 141
2 144 1 141
2 147 1 146
2 148 1 146
2 150 1 149
2 151 1 149
2 153 1 152
2 154 1 152
2 156 1 155
2 157 1 155
2 159 1 158
2 160 1 158
2 162 1 161
2 163 1 161
2 165 1 164
2 166 1 164
2 168 1 167
2 169 1 167
2 171 1 170
2 172 1 170
2 174 1 173
2 175 1 173
2 177 1 176
2 178 1 176
2 180 1 179
2 181 1 179
2 183 1 182
2 184 1 182
2 186 1 185
2 187 1 185
2 189 1 188
2 190 1 188
2 192 1 191
2 193 1 191
2 195 1 194
2 196 1 194
2 198 1 197
2 199 1 197
2 201 1 200
2 202 1 200
2 204 1 203
2 205 1 203
2 207 1 206
2 208 1 206
2 211 1 210
2 212 1 210
2 213 1 210
2 214 1 210
2 215 1 210
2 216 1 210
2 219 1 218
2 220 1 218
2 221 1 218
2 222 1 218
2 223 1 218
2 224 1 218
2 227 1 226
2 228 1 226
2 229 1 226
2 230 1 226
2 231 1 226
2 232 1 226
2 235 1 234
2 236 1 234
2 237 1 234
2 238 1 234
2 239 1 234
2 240 1 234
2 243 1 242
2 244 1 242
2 246 1 245
2 247 1 245
2 249 1 248
2 250 1 248
2 252 1 251
2 253 1 251
2 255 1 254
2 256 1 254
2 258 1 257
2 259 1 257
2 260 1 257
2 261 1 257
2 262 1 257
2 263 1 257
2 266 1 265
2 267 1 265
2 268 1 265
2 269 1 265
2 270 1 265
2 271 1 265
2 274 1 273
2 275 1 273
2 276 1 273
2 277 1 273
2 278 1 273
2 279 1 273
2 282 1 281
2 283 1 281
2 284 1 281
2 285 1 281
2 286 1 281
2 287 1 281
2 290 1 289
2 291 1 289
2 294 1 293
2 295 1 293
2 296 1 293
2 297 1 293
2 298 1 293
2 300 1 299
2 301 1 299
2 303 1 302
2 304 1 302
2 305 1 302
2 306 1 302
2 309 1 308
2 310 1 308
2 311 1 308
2 312 1 308
2 313 1 308
2 314 1 308
2 317 1 316
2 318 1 316
2 319 1 316
2 320 1 316
2 321 1 316
2 322 1 316
2 325 1 324
2 326 1 324
2 327 1 324
2 328 1 324
2 329 1 324
2 330 1 324
2 333 1 332
2 334 1 332
2 336 1 335
2 337 1 335
2 339 1 338
2 340 1 338
2 342 1 341
2 343 1 341
2 344 1 341
2 345 1 341
2 346 1 341
2 347 1 341
2 349 1 348
2 350 1 348
2 352 1 351
2 353 1 351
2 354 1 351
2 355 1 351
2 356 1 351
2 357 1 351
2 359 1 358
2 360 1 358
2 362 1 361
2 363 1 361
2 364 1 361
2 365 1 361
2 367 1 366
2 368 1 366
2 370 1 369
2 371 1 369
2 375 1 374
2 376 1 374
2 377 1 374
2 378 1 374
2 379 1 374
2 380 1 374
2 381 1 374
2 382 1 374
2 383 1 374
2 384 1 374
2 385 1 374
2 387 1 386
2 388 1 386
2 390 1 389
2 391 1 389
2 392 1 389
2 393 1 389
2 394 1 389
2 395 1 389
2 396 1 389
2 397 1 389
2 398 1 389
2 399 1 389
2 401 1 400
2 402 1 400
2 403 1 400
2 404 1 400
2 405 1 400
2 406 1 400
2 407 1 400
2 408 1 400
2 409 1 400
2 410 1 400
2 412 1 411
2 413 1 411
2 414 1 411
2 415 1 411
2 416 1 411
2 417 1 411
2 418 1 411
2 419 1 411
2 420 1 411
2 421 1 411
2 423 1 422
2 424 1 422
2 425 1 422
2 426 1 422
2 427 1 422
2 428 1 422
2 429 1 422
2 430 1 422
2 431 1 422
2 432 1 422
2 433 1 422
2 434 1 422
2 436 1 435
2 437 1 435
2 438 1 435
2 439 1 435
2 440 1 435
2 441 1 435
2 442 1 435
2 443 1 435
2 444 1 435
2 445 1 435
2 447 1 446
2 448 1 446
2 449 1 446
2 450 1 446
2 451 1 446
2 452 1 446
2 453 1 446
2 454 1 446
2 455 1 446
2 456 1 446
2 458 1 457
2 459 1 457
2 460 1 457
2 461 1 457
2 462 1 457
2 463 1 457
2 464 1 457
2 465 1 457
2 466 1 457
2 467 1 457
2 469 1 468
2 470 1 468
2 471 1 468
2 472 1 468
2 473 1 468
2 474 1 468
2 475 1 468
2 476 1 468
2 477 1 468
2 478 1 468
2 480 1 479
2 481 1 479
2 482 1 479
2 483 1 479
2 484 1 479
2 485 1 479
2 486 1 479
2 487 1 479
2 488 1 479
2 489 1 479
2 491 1 490
2 492 1 490
2 493 1 490
2 494 1 490
2 495 1 490
2 496 1 490
2 497 1 490
2 498 1 490
2 499 1 490
2 500 1 490
2 501 1 490
2 502 1 490
2 504 1 503
2 505 1 503
2 506 1 503
2 507 1 503
2 508 1 503
2 509 1 503
2 510 1 503
2 511 1 503
2 512 1 503
2 513 1 503
2 515 1 514
2 516 1 514
2 517 1 514
2 518 1 514
2 519 1 514
2 520 1 514
2 521 1 514
2 522 1 514
2 524 1 523
2 525 1 523
2 526 1 523
2 527 1 523
2 528 1 523
2 529 1 523
2 530 1 523
2 531 1 523
2 532 1 523
2 533 1 523
2 535 1 534
2 536 1 534
2 537 1 534
2 538 1 534
2 539 1 534
2 540 1 534
2 541 1 534
2 542 1 534
2 543 1 534
2 544 1 534
2 546 1 545
2 547 1 545
2 548 1 545
2 550 1 549
2 551 1 549
2 553 1 552
2 554 1 552
2 555 1 552
2 557 1 556
2 558 1 556
2 560 1 559
2 561 1 559
2 563 1 562
2 564 1 562
2 565 1 562
2 567 1 566
2 568 1 566
2 569 1 566
2 570 1 566
2 572 1 571
2 573 1 571
2 575 1 574
2 576 1 574
2 578 1 577
2 579 1 577
2 581 1 580
2 582 1 580
2 584 1 583
2 585 1 583
2 586 1 583
2 587 1 583
2 589 1 588
2 590 1 588
2 593 1 592
2 594 1 592
2 600 1 599
2 601 1 599
2 602 1 599
2 604 1 603
2 605 1 603
2 606 1 603
2 608 1 607
2 609 1 607
2 611 1 610
2 612 1 610
2 614 1 613
2 615 1 613
2 617 1 616
2 618 1 616
2 620 1 619
2 621 1 619
2 622 1 619
2 623 1 619
2 624 1 619
2 626 1 625
2 627 1 625
2 628 1 625
2 629 1 625
2 630 1 625
2 1068 1 1067
2 1069 1 1067
2 1070 1 1067
2 1071 1 1067
2 1072 1 1067
2 1073 1 1067
2 1074 1 1067
2 1075 1 1067
2 1076 1 1067
2 1077 1 1067
2 1078 1 1067
2 1079 1 1067
2 1081 1 1080
2 1082 1 1080
2 1083 1 1080
2 1084 1 1080
2 1085 1 1080
2 1086 1 1080
2 1087 1 1080
2 1088 1 1080
2 1089 1 1080
2 1090 1 1080
2 1091 1 1080
2 1093 1 1092
2 1094 1 1092
2 1095 1 1092
2 1096 1 1092
2 1097 1 1092
2 1098 1 1092
2 1099 1 1092
2 1100 1 1092
2 1101 1 1092
2 1102 1 1092
2 1103 1 1092
2 1105 1 1104
2 1106 1 1104
2 1107 1 1104
2 1108 1 1104
2 1109 1 1104
2 1110 1 1104
2 1111 1 1104
2 1112 1 1104
2 1113 1 1104
2 1114 1 1104
2 1115 1 1104
2 1116 1 1104
2 1158 1 1157
2 1159 1 1157
2 1160 1 1157
2 1162 1 1161
2 1163 1 1161
2 1164 1 1161
2 1165 1 1161
2 1166 1 1161
2 1167 1 1161
2 1168 1 1161
2 1169 1 1161
2 1170 1 1161
2 1171 1 1161
2 1172 1 1161
2 1174 1 1173
2 1175 1 1173
2 1176 1 1173
2 1177 1 1173
2 1178 1 1173
2 1179 1 1173
2 1180 1 1173
2 1181 1 1173
2 1182 1 1173
2 1183 1 1173
2 1184 1 1173
2 1186 1 1185
2 1187 1 1185
2 1188 1 1185
2 1189 1 1185
2 1190 1 1185
2 1191 1 1185
2 1192 1 1185
2 1193 1 1185
2 1194 1 1185
2 1195 1 1185
2 1196 1 1185
2 1198 1 1197
2 1199 1 1197
2 1200 1 1197
2 1201 1 1197
2 1202 1 1197
2 1203 1 1197
2 1204 1 1197
2 1205 1 1197
2 1206 1 1197
2 1207 1 1197
2 1208 1 1197
2 1210 1 1209
2 1211 1 1209
2 1212 1 1209
2 1214 1 1213
2 1215 1 1213
2 1217 1 1216
2 1218 1 1216
2 1220 1 1219
2 1221 1 1219
2 1222 1 1219
2 1224 1 1223
2 1225 1 1223
2 1226 1 1223
2 1227 1 1223
2 1228 1 1223
2 1229 1 1223
2 1230 1 1223
2 1231 1 1223
2 1232 1 1223
2 1233 1 1223
2 1234 1 1223
2 1236 1 1235
2 1237 1 1235
2 1238 1 1235
2 1239 1 1235
2 1240 1 1235
2 1241 1 1235
2 1242 1 1235
2 1243 1 1235
2 1244 1 1235
2 1245 1 1235
2 1246 1 1235
2 1248 1 1247
2 1249 1 1247
2 1250 1 1247
2 1251 1 1247
2 1252 1 1247
2 1253 1 1247
2 1254 1 1247
2 1255 1 1247
2 1256 1 1247
2 1257 1 1247
2 1258 1 1247
2 1260 1 1259
2 1261 1 1259
2 1262 1 1259
2 1263 1 1259
2 1264 1 1259
2 1265 1 1259
2 1266 1 1259
2 1267 1 1259
2 1268 1 1259
2 1269 1 1259
2 1270 1 1259
2 1272 1 1271
2 1273 1 1271
2 1274 1 1271
2 1275 1 1271
2 1276 1 1271
2 1277 1 1271
2 1278 1 1271
2 1279 1 1271
2 1281 1 1280
2 1282 1 1280
2 1283 1 1280
2 1284 1 1280
2 1285 1 1280
2 1286 1 1280
2 1287 1 1280
2 1288 1 1280
2 1289 1 1280
2 1290 1 1280
2 1291 1 1280
2 1293 1 1292
2 1294 1 1292
2 1295 1 1292
2 1296 1 1292
2 1297 1 1292
2 1298 1 1292
2 1299 1 1292
2 1300 1 1292
2 1301 1 1292
2 1302 1 1292
2 1304 1 1303
2 1305 1 1303
2 1306 1 1303
2 1307 1 1303
2 1308 1 1303
2 1309 1 1303
2 1310 1 1303
2 1311 1 1303
2 1312 1 1303
2 1313 1 1303
2 1314 1 1303
2 1316 1 1315
2 1317 1 1315
2 1318 1 1315
2 1319 1 1315
2 1320 1 1315
2 1321 1 1315
2 1322 1 1315
2 1323 1 1315
2 1324 1 1315
2 1325 1 1315
2 1326 1 1315
2 1328 1 1327
2 1329 1 1327
2 1330 1 1327
2 1331 1 1327
2 1332 1 1327
2 1333 1 1327
2 1334 1 1327
2 1335 1 1327
2 1336 1 1327
2 1337 1 1327
2 1338 1 1327
2 1340 1 1339
2 1341 1 1339
2 1342 1 1339
2 1343 1 1339
2 1344 1 1339
2 1345 1 1339
2 1346 1 1339
2 1347 1 1339
2 1348 1 1339
2 1349 1 1339
2 1350 1 1339
2 1352 1 1351
2 1353 1 1351
2 1354 1 1351
2 1355 1 1351
2 1356 1 1351
2 1357 1 1351
2 1358 1 1351
2 1359 1 1351
2 1360 1 1351
2 1361 1 1351
2 1362 1 1351
2 1364 1 1363
2 1365 1 1363
2 1366 1 1363
2 1367 1 1363
2 1368 1 1363
2 1369 1 1363
2 1370 1 1363
2 1371 1 1363
2 1372 1 1363
2 1373 1 1363
2 1374 1 1363
2 1376 1 1375
2 1377 1 1375
2 1379 1 1378
2 1380 1 1378
2 1382 1 1381
2 1383 1 1381
2 1385 1 1384
2 1386 1 1384
2 1388 1 1387
2 1389 1 1387
2 1391 1 1390
2 1392 1 1390
2 1394 1 1393
2 1395 1 1393
2 1397 1 1396
2 1398 1 1396
2 1416 1 1415
2 1417 1 1415
2 1419 1 1418
2 1420 1 1418
2 1422 1 1421
2 1423 1 1421
2 1425 1 1424
2 1426 1 1424
2 1428 1 1427
2 1429 1 1427
2 1431 1 1430
2 1432 1 1430
2 1434 1 1433
2 1435 1 1433
2 1437 1 1436
2 1438 1 1436
2 1456 1 1455
2 1457 1 1455
2 1458 1 1455
2 1459 1 1455
2 1460 1 1455
2 1461 1 1455
2 1463 1 1462
2 1464 1 1462
2 1465 1 1462
2 1466 1 1462
2 1467 1 1462
2 1468 1 1462
2 1470 1 1469
2 1471 1 1469
2 1472 1 1469
2 1473 1 1469
2 1474 1 1469
2 1476 1 1475
2 1477 1 1475
2 1478 1 1475
2 1480 1 1479
2 1481 1 1479
2 1483 1 1482
2 1484 1 1482
2 1485 1 1482
2 1486 1 1482
2 1487 1 1482
2 1488 1 1482
2 1489 1 1482
2 1490 1 1482
2 1491 1 1482
2 1493 1 1492
2 1494 1 1492
2 1496 1 1495
2 1497 1 1495
2 1499 1 1498
2 1500 1 1498
2 1502 1 1501
2 1503 1 1501
2 1505 1 1504
2 1506 1 1504
2 1508 1 1507
2 1509 1 1507
2 1511 1 1510
2 1512 1 1510
2 1514 1 1513
2 1515 1 1513
2 1517 1 1516
2 1518 1 1516
2 1520 1 1519
2 1521 1 1519
2 1523 1 1522
2 1524 1 1522
2 1526 1 1525
2 1527 1 1525
2 1543 1 1542
2 1544 1 1542
2 1546 1 1545
2 1547 1 1545
2 1549 1 1548
2 1550 1 1548
2 1552 1 1551
2 1553 1 1551
2 1555 1 1554
2 1556 1 1554
2 1558 1 1557
2 1559 1 1557
2 1561 1 1560
2 1562 1 1560
2 1564 1 1563
2 1565 1 1563
2 1567 1 1566
2 1568 1 1566
2 1569 1 1566
2 1570 1 1566
2 1571 1 1566
2 1572 1 1566
2 1574 1 1573
2 1575 1 1573
2 1576 1 1573
2 1577 1 1573
2 1578 1 1573
2 1579 1 1573
2 1581 1 1580
2 1582 1 1580
2 1584 1 1583
2 1585 1 1583
2 1586 1 1583
2 1587 1 1583
2 1589 1 1588
2 1590 1 1588
2 1591 1 1588
2 1592 1 1588
2 1593 1 1588
2 1595 1 1594
2 1596 1 1594
2 1598 1 1597
2 1599 1 1597
2 1601 1 1600
2 1602 1 1600
2 1604 1 1603
2 1605 1 1603
2 1607 1 1606
2 1608 1 1606
2 1610 1 1609
2 1611 1 1609
2 1613 1 1612
2 1614 1 1612
2 1616 1 1615
2 1617 1 1615
2 1619 1 1618
2 1620 1 1618
2 1622 1 1621
2 1623 1 1621
2 1625 1 1624
2 1626 1 1624
2 1628 1 1627
2 1629 1 1627
2 1631 1 1630
2 1632 1 1630
2 1634 1 1633
2 1635 1 1633
2 1637 1 1636
2 1638 1 1636
2 1640 1 1639
2 1641 1 1639
2 1643 1 1642
2 1644 1 1642
2 1646 1 1645
2 1647 1 1645
2 1649 1 1648
2 1650 1 1648
2 1652 1 1651
2 1653 1 1651
2 1655 1 1654
2 1656 1 1654
2 1658 1 1657
2 1659 1 1657
2 1661 1 1660
2 1662 1 1660
2 1664 1 1663
2 1665 1 1663
2 1666 1 1663
2 1667 1 1663
2 1668 1 1663
2 1669 1 1663
2 1670 1 1663
2 1671 1 1663
2 1672 1 1663
2 1673 1 1663
2 1674 1 1663
2 1676 1 1675
2 1677 1 1675
2 1678 1 1675
2 1679 1 1675
2 1680 1 1675
2 1681 1 1675
2 1682 1 1675
2 1683 1 1675
2 1684 1 1675
2 1686 1 1685
2 1687 1 1685
2 1688 1 1685
2 1689 1 1685
2 1690 1 1685
2 1691 1 1685
2 1692 1 1685
2 1693 1 1685
2 1694 1 1685
2 1695 1 1685
2 1696 1 1685
2 1698 1 1697
2 1699 1 1697
2 1700 1 1697
2 1701 1 1697
2 1702 1 1697
2 1703 1 1697
2 1704 1 1697
2 1705 1 1697
2 1706 1 1697
2 1707 1 1697
2 1708 1 1697
2 1710 1 1709
2 1711 1 1709
2 1712 1 1709
2 1713 1 1709
2 1714 1 1709
2 1715 1 1709
2 1716 1 1709
2 1717 1 1709
2 1718 1 1709
2 1719 1 1709
2 1720 1 1709
2 1722 1 1721
2 1723 1 1721
2 1724 1 1721
2 1725 1 1721
2 1726 1 1721
2 1728 1 1727
2 1729 1 1727
2 1730 1 1727
2 1732 1 1731
2 1733 1 1731
2 1734 1 1731
2 1735 1 1731
2 1736 1 1731
2 1737 1 1731
2 1738 1 1731
2 1739 1 1731
2 1740 1 1731
2 1741 1 1731
2 1742 1 1731
2 1744 1 1743
2 1745 1 1743
2 1746 1 1743
2 1747 1 1743
2 1748 1 1743
2 1749 1 1743
2 1750 1 1743
2 1751 1 1743
2 1752 1 1743
2 1753 1 1743
2 1754 1 1743
2 1756 1 1755
2 1757 1 1755
2 1759 1 1758
2 1760 1 1758
2 1762 1 1761
2 1763 1 1761
2 1764 1 1761
2 1765 1 1761
2 1766 1 1761
2 1767 1 1761
2 1768 1 1761
2 1770 1 1769
2 1771 1 1769
2 1772 1 1769
2 1773 1 1769
2 1774 1 1769
2 1775 1 1769
2 1776 1 1769
2 1778 1 1777
2 1779 1 1777
2 1780 1 1777
2 1781 1 1777
2 1782 1 1777
2 1783 1 1777
2 1784 1 1777
2 1786 1 1785
2 1787 1 1785
2 1788 1 1785
2 1789 1 1785
2 1790 1 1785
2 1791 1 1785
2 1792 1 1785
2 1794 1 1793
2 1795 1 1793
2 1796 1 1793
2 1797 1 1793
2 1798 1 1793
2 1799 1 1793
2 1801 1 1800
2 1802 1 1800
2 1803 1 1800
2 1804 1 1800
2 1805 1 1800
2 1806 1 1800
2 1808 1 1807
2 1809 1 1807
2 1810 1 1807
2 1811 1 1807
2 1812 1 1807
2 1813 1 1807
2 1815 1 1814
2 1816 1 1814
2 1817 1 1814
2 1818 1 1814
2 1819 1 1814
2 1820 1 1814
2 1822 1 1821
2 1823 1 1821
2 1825 1 1824
2 1826 1 1824
2 1828 1 1827
2 1829 1 1827
2 1831 1 1830
2 1832 1 1830
2 1834 1 1833
2 1835 1 1833
2 1837 1 1836
2 1838 1 1836
2 1840 1 1839
2 1841 1 1839
2 1843 1 1842
2 1844 1 1842
2 1846 1 1845
2 1847 1 1845
2 1849 1 1848
2 1850 1 1848
2 1852 1 1851
2 1853 1 1851
2 1855 1 1854
2 1856 1 1854
2 1858 1 1857
2 1859 1 1857
2 1861 1 1860
2 1862 1 1860
2 1864 1 1863
2 1865 1 1863
2 1867 1 1866
2 1868 1 1866
2 1870 1 1869
2 1871 1 1869
2 1873 1 1872
2 1874 1 1872
2 1876 1 1875
2 1877 1 1875
2 1879 1 1878
2 1880 1 1878
2 1882 1 1881
2 1883 1 1881
2 1885 1 1884
2 1886 1 1884
2 1888 1 1887
2 1889 1 1887
2 1891 1 1890
2 1892 1 1890
2 1894 1 1893
2 1895 1 1893
2 1897 1 1896
2 1898 1 1896
2 1900 1 1899
2 1901 1 1899
2 1903 1 1902
2 1904 1 1902
2 1906 1 1905
2 1907 1 1905
2 1909 1 1908
2 1910 1 1908
2 1912 1 1911
2 1913 1 1911
2 1915 1 1914
2 1916 1 1914
2 1918 1 1917
2 1919 1 1917
2 1921 1 1920
2 1922 1 1920
2 1924 1 1923
2 1925 1 1923
2 1927 1 1926
2 1928 1 1926
2 1930 1 1929
2 1931 1 1929
2 1933 1 1932
2 1934 1 1932
2 1936 1 1935
2 1937 1 1935
2 1939 1 1938
2 1940 1 1938
2 1942 1 1941
2 1943 1 1941
2 1945 1 1944
2 1946 1 1944
2 1948 1 1947
2 1949 1 1947
2 1951 1 1950
2 1952 1 1950
2 1954 1 1953
2 1955 1 1953
2 1957 1 1956
2 1958 1 1956
2 1960 1 1959
2 1961 1 1959
2 1963 1 1962
2 1964 1 1962
2 1966 1 1965
2 1967 1 1965
2 1969 1 1968
2 1970 1 1968
2 2648 1 2647
2 2649 1 2647
2 2650 1 2647
2 2651 1 2647
2 2652 1 2647
2 2654 1 2653
2 2655 1 2653
2 2656 1 2653
2 2657 1 2653
2 2658 1 2653
2 2659 1 2653
2 2660 1 2653
2 2661 1 2653
2 2662 1 2653
2 2663 1 2653
2 2665 1 2664
2 2666 1 2664
2 2667 1 2664
2 2668 1 2664
2 2669 1 2664
2 2670 1 2664
2 2671 1 2664
2 2672 1 2664
2 2673 1 2664
2 2674 1 2664
2 2676 1 2675
2 2677 1 2675
2 2678 1 2675
2 2679 1 2675
2 2680 1 2675
2 2682 1 2681
2 2683 1 2681
2 2684 1 2681
2 2685 1 2681
2 2686 1 2681
2 2687 1 2681
2 2688 1 2681
2 2689 1 2681
2 2690 1 2681
2 2691 1 2681
2 2693 1 2692
2 2694 1 2692
2 2695 1 2692
2 2696 1 2692
2 2697 1 2692
2 2698 1 2692
2 2699 1 2692
2 2700 1 2692
2 2701 1 2692
2 2702 1 2692
2 2705 1 2704
2 2706 1 2704
2 2707 1 2704
2 2708 1 2704
2 2723 1 2722
2 2724 1 2722
2 2725 1 2722
2 2726 1 2722
2 2727 1 2722
2 2729 1 2728
2 2730 1 2728
2 2731 1 2728
2 2732 1 2728
2 2733 1 2728
2 2734 1 2728
2 2735 1 2728
2 2736 1 2728
2 2737 1 2728
2 2738 1 2728
2 2740 1 2739
2 2741 1 2739
2 2742 1 2739
2 2743 1 2739
2 2744 1 2739
2 2745 1 2739
2 2746 1 2739
2 2747 1 2739
2 2748 1 2739
2 2749 1 2739
2 2751 1 2750
2 2752 1 2750
2 2753 1 2750
2 2754 1 2750
2 2755 1 2750
2 2757 1 2756
2 2758 1 2756
2 2759 1 2756
2 2760 1 2756
2 2761 1 2756
2 2762 1 2756
2 2763 1 2756
2 2764 1 2756
2 2765 1 2756
2 2766 1 2756
2 2768 1 2767
2 2769 1 2767
2 2770 1 2767
2 2771 1 2767
2 2772 1 2767
2 2773 1 2767
2 2774 1 2767
2 2775 1 2767
2 2776 1 2767
2 2777 1 2767
2 2780 1 2779
2 2781 1 2779
2 2782 1 2779
2 2783 1 2779
2 2784 1 2779
2 2785 1 2779
2 2786 1 2779
2 2787 1 2779
2 2788 1 2779
2 2789 1 2779
2 2791 1 2790
2 2792 1 2790
2 2793 1 2790
2 2794 1 2790
2 2795 1 2790
2 2796 1 2790
2 2797 1 2790
2 2798 1 2790
2 2799 1 2790
2 2800 1 2790
2 2802 1 2801
2 2803 1 2801
2 2804 1 2801
2 2805 1 2801
2 2806 1 2801
2 2807 1 2801
2 2808 1 2801
2 2809 1 2801
2 2810 1 2801
2 2811 1 2801
2 2813 1 2812
2 2814 1 2812
2 2815 1 2812
2 2816 1 2812
2 2817 1 2812
2 2818 1 2812
2 2819 1 2812
2 2820 1 2812
2 2821 1 2812
2 2822 1 2812
2 2856 1 2855
2 2857 1 2855
2 2858 1 2855
2 2859 1 2855
2 2860 1 2855
2 2862 1 2861
2 2863 1 2861
2 2864 1 2861
2 2865 1 2861
2 2866 1 2861
2 2878 1 2877
2 2879 1 2877
2 2880 1 2877
2 2881 1 2877
2 2883 1 2882
2 2884 1 2882
2 2885 1 2882
2 2886 1 2882
2 2887 1 2882
2 2888 1 2882
2 2889 1 2882
2 2890 1 2882
2 2892 1 2891
2 2893 1 2891
2 2894 1 2891
2 2895 1 2891
2 2896 1 2891
2 2897 1 2891
2 2898 1 2891
2 2899 1 2891
2 2900 1 2891
2 2943 1 2942
2 2944 1 2942
2 2945 1 2942
2 2946 1 2942
2 2947 1 2942
2 2949 1 2948
2 2950 1 2948
2 2951 1 2948
2 2952 1 2948
2 2953 1 2948
2 2965 1 2964
2 2966 1 2964
2 2967 1 2964
2 2968 1 2964
2 3001 1 3000
2 3002 1 3000
2 3004 1 3003
2 3005 1 3003
2 3008 1 3007
2 3009 1 3007
2 3011 1 3010
2 3012 1 3010
2 3036 1 3035
2 3037 1 3035
2 3039 1 3038
2 3040 1 3038
2 3042 1 3041
2 3043 1 3041
2 3044 1 3041
2 3045 1 3041
2 3046 1 3041
2 3047 1 3041
2 3048 1 3041
2 3049 1 3041
2 3050 1 3041
2 3051 1 3041
2 3053 1 3052
2 3054 1 3052
2 3055 1 3052
2 3056 1 3052
2 3057 1 3052
2 3058 1 3052
2 3059 1 3052
2 3060 1 3052
2 3061 1 3052
2 3062 1 3052
2 3064 1 3063
2 3065 1 3063
2 3066 1 3063
2 3067 1 3063
2 3069 1 3068
2 3070 1 3068
2 3076 1 3075
2 3077 1 3075
2 3078 1 3075
2 3079 1 3075
2 3080 1 3075
2 3081 1 3075
2 3082 1 3075
2 3083 1 3075
2 3084 1 3075
2 3085 1 3075
2 3087 1 3086
2 3088 1 3086
2 3089 1 3086
2 3090 1 3086
2 3091 1 3086
2 3092 1 3086
2 3093 1 3086
2 3094 1 3086
2 3095 1 3086
2 3096 1 3086
2 3098 1 3097
2 3099 1 3097
2 3100 1 3097
2 3101 1 3097
2 3102 1 3097
2 3103 1 3097
2 3104 1 3097
2 3105 1 3097
2 3106 1 3097
2 3107 1 3097
2 3109 1 3108
2 3110 1 3108
2 3111 1 3108
2 3112 1 3108
2 3113 1 3108
2 3114 1 3108
2 3115 1 3108
2 3116 1 3108
2 3117 1 3108
2 3118 1 3108
2 3120 1 3119
2 3121 1 3119
2 3122 1 3119
2 3123 1 3119
2 3124 1 3119
2 3125 1 3119
2 3126 1 3119
2 3127 1 3119
2 3128 1 3119
2 3129 1 3119
2 3131 1 3130
2 3132 1 3130
2 3133 1 3130
2 3134 1 3130
2 3135 1 3130
2 3136 1 3130
2 3137 1 3130
2 3138 1 3130
2 3139 1 3130
2 3140 1 3130
2 3148 1 3147
2 3149 1 3147
2 3150 1 3147
2 3151 1 3147
2 3152 1 3147
2 3153 1 3147
2 3154 1 3147
2 3155 1 3147
2 3156 1 3147
2 3157 1 3147
2 3159 1 3158
2 3160 1 3158
2 3161 1 3158
2 3162 1 3158
2 3163 1 3158
2 3164 1 3158
2 3165 1 3158
2 3166 1 3158
2 3167 1 3158
2 3168 1 3158
2 3170 1 3169
2 3171 1 3169
2 3172 1 3169
2 3173 1 3169
2 3174 1 3169
2 3175 1 3169
2 3176 1 3169
2 3177 1 3169
2 3178 1 3169
2 3179 1 3169
2 3181 1 3180
2 3182 1 3180
2 3183 1 3180
2 3184 1 3180
2 3185 1 3180
2 3186 1 3180
2 3187 1 3180
2 3188 1 3180
2 3189 1 3180
2 3190 1 3180
2 3192 1 3191
2 3193 1 3191
2 3201 1 3200
2 3202 1 3200
2 3457 1 3456
2 3458 1 3456
2 3692 1 3691
2 3693 1 3691
2 3694 1 3691
2 3695 1 3691
2 3696 1 3691
2 3697 1 3691
2 3698 1 3691
2 3699 1 3691
2 3706 1 3705
2 3707 1 3705
2 3733 1 3732
2 3734 1 3732
2 3735 1 3732
2 3736 1 3732
2 3737 1 3732
2 3772 1 3771
2 3773 1 3771
2 3774 1 3771
2 3776 1 3775
2 3777 1 3775
2 3778 1 3775
2 3790 1 3789
2 3791 1 3789
2 3792 1 3789
2 3794 1 3793
2 3795 1 3793
2 3796 1 3793
2 3798 1 3797
2 3799 1 3797
2 3811 1 3810
2 3812 1 3810
2 3814 1 3813
2 3815 1 3813
2 3817 1 3816
2 3818 1 3816
2 3820 1 3819
2 3821 1 3819
2 3825 1 3824
2 3826 1 3824
2 3843 1 3842
2 3844 1 3842
2 3845 1 3842
2 3846 1 3842
2 3847 1 3842
2 3848 1 3842
2 3850 1 3849
2 3851 1 3849
2 3852 1 3849
2 3853 1 3849
2 3854 1 3849
2 3856 1 3855
2 3857 1 3855
2 3858 1 3855
2 3859 1 3855
2 3860 1 3855
2 3862 1 3861
2 3863 1 3861
2 3864 1 3861
2 3865 1 3861
2 3866 1 3861
2 3868 1 3867
2 3869 1 3867
2 3870 1 3867
2 3871 1 3867
2 3872 1 3867
2 3874 1 3873
2 3875 1 3873
2 3876 1 3873
2 3877 1 3873
2 3878 1 3873
2 3879 1 3873
2 3880 1 3873
2 3882 1 3881
2 3883 1 3881
2 3884 1 3881
2 3885 1 3881
2 3886 1 3881
2 3888 1 3887
2 3889 1 3887
2 3890 1 3887
2 3891 1 3887
2 3892 1 3887
2 3894 1 3893
2 3895 1 3893
2 3896 1 3893
2 3897 1 3893
2 3898 1 3893
2 3912 1 3911
2 3913 1 3911
2 3922 1 3921
2 3923 1 3921
2 3924 1 3921
2 3925 1 3921
2 3926 1 3921
2 3928 1 3927
2 3929 1 3927
2 3930 1 3927
2 3931 1 3927
2 3932 1 3927
2 3934 1 3933
2 3935 1 3933
2 3936 1 3933
2 3937 1 3933
2 3938 1 3933
2 3943 1 3942
2 3944 1 3942
2 3945 1 3942
2 3946 1 3942
2 3947 1 3942
2 3949 1 3948
2 3950 1 3948
2 3951 1 3948
2 3952 1 3948
2 3953 1 3948
2 3954 1 3948
2 3955 1 3948
2 3957 1 3956
2 3958 1 3956
2 3959 1 3956
2 3960 1 3956
2 3961 1 3956
2 3963 1 3962
2 3964 1 3962
2 3965 1 3962
2 3966 1 3962
2 3967 1 3962
2 3969 1 3968
2 3970 1 3968
2 3971 1 3968
2 3972 1 3968
2 3973 1 3968
2 3974 1 3968
2 3985 1 3984
2 3986 1 3984
2 4009 1 4008
2 4010 1 4008
2 4012 1 4011
2 4013 1 4011
2 4022 1 4021
2 4023 1 4021
2 4068 1 4067
2 4069 1 4067
2 4081 1 4080
2 4082 1 4080
2 4083 1 4080
2 4089 1 4088
2 4090 1 4088
2 4092 1 4091
2 4093 1 4091
2 4095 1 4094
2 4096 1 4094
2 4098 1 4097
2 4099 1 4097
2 4101 1 4100
2 4102 1 4100
2 4104 1 4103
2 4105 1 4103
2 4107 1 4106
2 4108 1 4106
2 4110 1 4109
2 4111 1 4109
2 4145 1 4144
2 4146 1 4144
2 4148 1 4147
2 4149 1 4147
2 4151 1 4150
2 4152 1 4150
2 4154 1 4153
2 4155 1 4153
2 4157 1 4156
2 4158 1 4156
2 4160 1 4159
2 4161 1 4159
2 4189 1 4188
2 4190 1 4188
2 4192 1 4191
2 4193 1 4191
2 4201 1 4200
2 4202 1 4200
2 4204 1 4203
2 4205 1 4203
2 4207 1 4206
2 4208 1 4206
2 4210 1 4209
2 4211 1 4209
2 4213 1 4212
2 4214 1 4212
2 4216 1 4215
2 4217 1 4215
2 4220 1 4219
2 4221 1 4219
2 4226 1 4225
2 4227 1 4225
2 4229 1 4228
2 4230 1 4228
2 4232 1 4231
2 4233 1 4231
2 4235 1 4234
2 4236 1 4234
2 4238 1 4237
2 4239 1 4237
2 4241 1 4240
2 4242 1 4240
2 4244 1 4243
2 4245 1 4243
2 4247 1 4246
2 4248 1 4246
2 4250 1 4249
2 4251 1 4249
2 4253 1 4252
2 4254 1 4252
2 4256 1 4255
2 4257 1 4255
2 4259 1 4258
2 4260 1 4258
2 4265 1 4264
2 4266 1 4264
2 4281 1 4280
2 4282 1 4280
2 4283 1 4280
2 4285 1 4284
2 4286 1 4284
2 4287 1 4284
2 4288 1 4284
2 4289 1 4284
2 4291 1 4290
2 4292 1 4290
2 4293 1 4290
2 4294 1 4290
2 4295 1 4290
2 4296 1 4290
2 4299 1 4298
2 4300 1 4298
2 4302 1 4301
2 4303 1 4301
2 4304 1 4301
2 4306 1 4305
2 4307 1 4305
2 4308 1 4305
2 4309 1 4305
2 4311 1 4310
2 4312 1 4310
2 4313 1 4310
2 4314 1 4310
2 4315 1 4310
2 4317 1 4316
2 4318 1 4316
2 4319 1 4316
2 4321 1 4320
2 4322 1 4320
2 4323 1 4320
2 4324 1 4320
2 4326 1 4325
2 4327 1 4325
2 4328 1 4325
2 4329 1 4325
2 4330 1 4325
2 4333 1 4332
2 4334 1 4332
2 4335 1 4332
2 4337 1 4336
2 4338 1 4336
2 4339 1 4336
2 4340 1 4336
2 4341 1 4336
2 4343 1 4342
2 4344 1 4342
2 4345 1 4342
2 4346 1 4342
2 4347 1 4342
2 4348 1 4342
2 4350 1 4349
2 4351 1 4349
2 4352 1 4349
2 4353 1 4349
2 4354 1 4349
2 4355 1 4349
2 4356 1 4349
2 4358 1 4357
2 4359 1 4357
2 4360 1 4357
2 4361 1 4357
2 4362 1 4357
2 4363 1 4357
2 4365 1 4364
2 4366 1 4364
2 4367 1 4364
2 4368 1 4364
2 4369 1 4364
2 4370 1 4364
2 4371 1 4364
2 4372 1 4364
2 4373 1 4364
2 4374 1 4364
2 4376 1 4375
2 4377 1 4375
2 4378 1 4375
2 4380 1 4379
2 4381 1 4379
2 4382 1 4379
2 4383 1 4379
2 4384 1 4379
2 4386 1 4385
2 4387 1 4385
2 4388 1 4385
2 4389 1 4385
2 4390 1 4385
2 4391 1 4385
2 4397 1 4396
2 4398 1 4396
2 4399 1 4396
2 4401 1 4400
2 4402 1 4400
2 4403 1 4400
2 4404 1 4400
2 4406 1 4405
2 4407 1 4405
2 4408 1 4405
2 4409 1 4405
2 4410 1 4405
2 4411 1 4405
2 4413 1 4412
2 4414 1 4412
2 4415 1 4412
2 4416 1 4412
2 4417 1 4412
2 4419 1 4418
2 4420 1 4418
2 4421 1 4418
2 4422 1 4418
2 4423 1 4418
2 4424 1 4418
2 4426 1 4425
2 4427 1 4425
2 4428 1 4425
2 4429 1 4425
2 4430 1 4425
2 4431 1 4425
2 4432 1 4425
2 4433 1 4425
2 4434 1 4425
2 4435 1 4425
2 4437 1 4436
2 4438 1 4436
2 4439 1 4436
2 4441 1 4440
2 4442 1 4440
2 4443 1 4440
2 4444 1 4440
2 4446 1 4445
2 4447 1 4445
2 4448 1 4445
2 4449 1 4445
2 4450 1 4445
2 4457 1 4456
2 4458 1 4456
2 4459 1 4456
2 4460 1 4456
2 4461 1 4456
2 4463 1 4462
2 4464 1 4462
2 4465 1 4462
2 4466 1 4462
2 4467 1 4462
2 4468 1 4462
2 4470 1 4469
2 4471 1 4469
2 4472 1 4469
2 4473 1 4469
2 4474 1 4469
2 4475 1 4469
2 4476 1 4469
2 4478 1 4477
2 4479 1 4477
2 4480 1 4477
2 4481 1 4477
2 4482 1 4477
2 4483 1 4477
2 4513 1 4512
2 4514 1 4512
2 4525 1 4524
2 4526 1 4524
2 4527 1 4524
2 4533 1 4532
2 4534 1 4532
2 4535 1 4532
2 4549 1 4548
2 4550 1 4548
2 4552 1 4551
2 4553 1 4551
2 4555 1 4554
2 4556 1 4554
2 4558 1 4557
2 4559 1 4557
2 4561 1 4560
2 4562 1 4560
2 4564 1 4563
2 4565 1 4563
2 4567 1 4566
2 4568 1 4566
2 4570 1 4569
2 4571 1 4569
2 4573 1 4572
2 4574 1 4572
2 4576 1 4575
2 4577 1 4575
2 4579 1 4578
2 4580 1 4578
2 4582 1 4581
2 4583 1 4581
2 4585 1 4584
2 4586 1 4584
2 4588 1 4587
2 4589 1 4587
2 4591 1 4590
2 4592 1 4590
2 4594 1 4593
2 4595 1 4593
2 4597 1 4596
2 4598 1 4596
2 4600 1 4599
2 4601 1 4599
2 4603 1 4602
2 4604 1 4602
2 4606 1 4605
2 4607 1 4605
2 4609 1 4608
2 4610 1 4608
2 4612 1 4611
2 4613 1 4611
2 4615 1 4614
2 4616 1 4614
2 4618 1 4617
2 4619 1 4617
2 4622 1 4621
2 4623 1 4621
2 4625 1 4624
2 4626 1 4624
2 4628 1 4627
2 4629 1 4627
2 4631 1 4630
2 4632 1 4630
2 4634 1 4633
2 4635 1 4633
2 4638 1 4637
2 4639 1 4637
2 4641 1 4640
2 4642 1 4640
2 4644 1 4643
2 4645 1 4643
2 4647 1 4646
2 4648 1 4646
2 4650 1 4649
2 4651 1 4649
2 4653 1 4652
2 4654 1 4652
2 4656 1 4655
2 4657 1 4655
2 4659 1 4658
2 4660 1 4658
2 4663 1 4662
2 4664 1 4662
2 4666 1 4665
2 4667 1 4665
2 4669 1 4668
2 4670 1 4668
2 4672 1 4671
2 4673 1 4671
2 4675 1 4674
2 4676 1 4674
2 4678 1 4677
2 4679 1 4677
2 4681 1 4680
2 4682 1 4680
2 4684 1 4683
2 4685 1 4683
2 4687 1 4686
2 4688 1 4686
2 4690 1 4689
2 4691 1 4689
2 4693 1 4692
2 4694 1 4692
2 4696 1 4695
2 4697 1 4695
2 4699 1 4698
2 4700 1 4698
2 4940 1 4939
2 4941 1 4939
2 5050 1 5049
2 5051 1 5049
2 5151 1 5150
2 5152 1 5150
2 5158 1 5157
2 5159 1 5157
2 5167 1 5166
2 5168 1 5166
2 5170 1 5169
2 5171 1 5169
2 5174 1 5173
2 5175 1 5173
2 5178 1 5177
2 5179 1 5177
2 5181 1 5180
2 5182 1 5180
2 5184 1 5183
2 5185 1 5183
2 5187 1 5186
2 5188 1 5186
2 5190 1 5189
2 5191 1 5189
2 5193 1 5192
2 5194 1 5192
2 5196 1 5195
2 5197 1 5195
2 5200 1 5199
2 5201 1 5199
2 5203 1 5202
2 5204 1 5202
2 5206 1 5205
2 5207 1 5205
2 5209 1 5208
2 5210 1 5208
2 5212 1 5211
2 5213 1 5211
2 5215 1 5214
2 5216 1 5214
2 5218 1 5217
2 5219 1 5217
2 5221 1 5220
2 5222 1 5220
2 5237 1 5236
2 5238 1 5236
2 5265 1 5264
2 5266 1 5264
2 5267 1 5264
2 5268 1 5264
2 5269 1 5264
2 5270 1 5264
2 5271 1 5264
2 5272 1 5264
2 5273 1 5264
2 5285 1 5284
2 5286 1 5284
2 5287 1 5284
2 5288 1 5284
2 5289 1 5284
2 5290 1 5284
2 5291 1 5284
2 5292 1 5284
2 5293 1 5284
2 5294 1 5284
2 5295 1 5284
2 5296 1 5284
2 5297 1 5284
2 5316 1 5315
2 5317 1 5315
2 5318 1 5315
2 5320 1 5319
2 5321 1 5319
2 5325 1 5324
2 5326 1 5324
2 5327 1 5324
2 5329 1 5328
2 5330 1 5328
2 5347 1 5346
2 5348 1 5346
2 5372 1 5371
2 5373 1 5371
2 5375 1 5374
2 5376 1 5374
2 5378 1 5377
2 5379 1 5377
2 5383 1 5382
2 5384 1 5382
2 5386 1 5385
2 5387 1 5385
2 5390 1 5389
2 5391 1 5389
2 5392 1 5389
2 5393 1 5389
2 5394 1 5389
2 5395 1 5389
2 5397 1 5396
2 5398 1 5396
2 5399 1 5396
2 5400 1 5396
2 5401 1 5396
2 5402 1 5396
2 5403 1 5396
2 5404 1 5396
2 5405 1 5396
2 5406 1 5396
2 5408 1 5407
2 5409 1 5407
2 5410 1 5407
2 5411 1 5407
2 5412 1 5407
2 5413 1 5407
2 5414 1 5407
2 5415 1 5407
2 5416 1 5407
2 5417 1 5407
2 5419 1 5418
2 5420 1 5418
2 5421 1 5418
2 5422 1 5418
2 5423 1 5418
2 5425 1 5424
2 5426 1 5424
2 5427 1 5424
2 5428 1 5424
2 5429 1 5424
2 5430 1 5424
2 5432 1 5431
2 5433 1 5431
2 5434 1 5431
2 5435 1 5431
2 5436 1 5431
2 5437 1 5431
2 5438 1 5431
2 5439 1 5431
2 5440 1 5431
2 5442 1 5441
2 5443 1 5441
2 5444 1 5441
2 5445 1 5441
2 5446 1 5441
2 5447 1 5441
2 5448 1 5441
2 5449 1 5441
2 5450 1 5441
2 5451 1 5441
2 5453 1 5452
2 5454 1 5452
2 5455 1 5452
2 5456 1 5452
2 5457 1 5452
2 5458 1 5452
2 5459 1 5452
2 5460 1 5452
2 5461 1 5452
2 5463 1 5462
2 5464 1 5462
2 5465 1 5462
2 5466 1 5462
2 5467 1 5462
2 5468 1 5462
2 5471 1 5470
2 5472 1 5470
2 5473 1 5470
2 5474 1 5470
2 5475 1 5470
2 5476 1 5470
2 5478 1 5477
2 5479 1 5477
2 5480 1 5477
2 5481 1 5477
2 5482 1 5477
2 5483 1 5477
2 5484 1 5477
2 5485 1 5477
2 5486 1 5477
2 5487 1 5477
2 5489 1 5488
2 5490 1 5488
2 5491 1 5488
2 5492 1 5488
2 5493 1 5488
2 5494 1 5488
2 5495 1 5488
2 5496 1 5488
2 5497 1 5488
2 5499 1 5498
2 5500 1 5498
2 5501 1 5498
2 5502 1 5498
2 5503 1 5498
2 5504 1 5498
2 5505 1 5498
2 5507 1 5506
2 5508 1 5506
2 5509 1 5506
2 5510 1 5506
2 5511 1 5506
2 5512 1 5506
2 5513 1 5506
2 5514 1 5506
2 5515 1 5506
2 5516 1 5506
2 5517 1 5506
2 5518 1 5506
2 5519 1 5506
2 5521 1 5520
2 5522 1 5520
2 5523 1 5520
2 5524 1 5520
2 5525 1 5520
2 5526 1 5520
2 5527 1 5520
2 5528 1 5520
2 5529 1 5520
2 5530 1 5520
2 5531 1 5520
2 5532 1 5520
2 5533 1 5520
2 5534 1 5520
2 5535 1 5520
2 5537 1 5536
2 5538 1 5536
2 5539 1 5536
2 5540 1 5536
2 5541 1 5536
2 5542 1 5536
2 5543 1 5536
2 5544 1 5536
2 5545 1 5536
2 5546 1 5536
2 5547 1 5536
2 5548 1 5536
2 5550 1 5549
2 5551 1 5549
2 5552 1 5549
2 5553 1 5549
2 5554 1 5549
2 5556 1 5555
2 5557 1 5555
2 5558 1 5555
2 5559 1 5555
2 5560 1 5555
2 5561 1 5555
2 5563 1 5562
2 5564 1 5562
2 5565 1 5562
2 5566 1 5562
2 5567 1 5562
2 5568 1 5562
2 5569 1 5562
2 5570 1 5562
2 5571 1 5562
2 5572 1 5562
2 5574 1 5573
2 5575 1 5573
2 5576 1 5573
2 5577 1 5573
2 5578 1 5573
2 5580 1 5579
2 5581 1 5579
2 5582 1 5579
2 5583 1 5579
2 5584 1 5579
2 5585 1 5579
2 5596 1 5595
2 5597 1 5595
2 5598 1 5595
2 5599 1 5595
2 5600 1 5595
2 5601 1 5595
2 5602 1 5595
2 5603 1 5595
2 5604 1 5595
2 5605 1 5595
2 5607 1 5606
2 5608 1 5606
2 5609 1 5606
2 5610 1 5606
2 5611 1 5606
2 5612 1 5606
2 5613 1 5606
2 5614 1 5606
2 5615 1 5606
2 5625 1 5624
2 5626 1 5624
2 5627 1 5624
2 5628 1 5624
2 5629 1 5624
2 5630 1 5624
2 5631 1 5624
2 5632 1 5624
2 5633 1 5624
2 5635 1 5634
2 5636 1 5634
2 5637 1 5634
2 5638 1 5634
2 5639 1 5634
2 5640 1 5634
2 5641 1 5634
2 5656 1 5655
2 5657 1 5655
2 5658 1 5655
2 5659 1 5655
2 5660 1 5655
2 5661 1 5655
2 5662 1 5655
2 5663 1 5655
2 5664 1 5655
2 5665 1 5655
2 5666 1 5655
2 5667 1 5655
2 5668 1 5655
2 5669 1 5655
2 5670 1 5655
2 5672 1 5671
2 5673 1 5671
2 5674 1 5671
2 5675 1 5671
2 5676 1 5671
2 5677 1 5671
2 5678 1 5671
2 5679 1 5671
2 5680 1 5671
2 5681 1 5671
2 5682 1 5671
2 5683 1 5671
2 5685 1 5684
2 5686 1 5684
2 5687 1 5684
2 5688 1 5684
2 5689 1 5684
2 5693 1 5692
2 5694 1 5692
2 5695 1 5692
2 5697 1 5696
2 5698 1 5696
2 5699 1 5696
2 5701 1 5700
2 5702 1 5700
2 5704 1 5703
2 5705 1 5703
2 5706 1 5703
2 5708 1 5707
2 5709 1 5707
2 5710 1 5707
2 5712 1 5711
2 5713 1 5711
2 5737 1 5736
2 5738 1 5736
2 5740 1 5739
2 5741 1 5739
2 5743 1 5742
2 5744 1 5742
2 5746 1 5745
2 5747 1 5745
2 5757 1 5756
2 5758 1 5756
2 6026 1 6025
2 6027 1 6025
2 6029 1 6028
2 6030 1 6028
2 6032 1 6031
2 6033 1 6031
2 6035 1 6034
2 6036 1 6034
2 6038 1 6037
2 6039 1 6037
2 6041 1 6040
2 6042 1 6040
2 6046 1 6045
2 6047 1 6045
2 6049 1 6048
2 6050 1 6048
2 6052 1 6051
2 6053 1 6051
2 6055 1 6054
2 6056 1 6054
2 6081 1 6080
2 6082 1 6080
2 6092 1 6091
2 6093 1 6091
2 6109 1 6108
2 6110 1 6108
2 6118 1 6117
2 6119 1 6117
2 6141 1 6140
2 6142 1 6140
2 6150 1 6149
2 6151 1 6149
2 6165 1 6164
2 6166 1 6164
2 6169 1 6168
2 6170 1 6168
2 6176 1 6175
2 6177 1 6175
2 6198 1 6197
2 6199 1 6197
2 6201 1 6200
2 6202 1 6200
2 6204 1 6203
2 6205 1 6203
2 6207 1 6206
2 6208 1 6206
2 6210 1 6209
2 6211 1 6209
2 6213 1 6212
2 6214 1 6212
2 6216 1 6215
2 6217 1 6215
2 6219 1 6218
2 6220 1 6218
2 6239 1 6238
2 6240 1 6238
2 6242 1 6241
2 6243 1 6241
2 6245 1 6244
2 6246 1 6244
2 6248 1 6247
2 6249 1 6247
2 6251 1 6250
2 6252 1 6250
2 6254 1 6253
2 6255 1 6253
2 6257 1 6256
2 6258 1 6256
2 6260 1 6259
2 6261 1 6259
2 6263 1 6262
2 6264 1 6262
2 6266 1 6265
2 6267 1 6265
2 6269 1 6268
2 6270 1 6268
2 6272 1 6271
2 6273 1 6271
2 6275 1 6274
2 6276 1 6274
2 6278 1 6277
2 6279 1 6277
2 6281 1 6280
2 6282 1 6280
2 6284 1 6283
2 6285 1 6283
2 6287 1 6286
2 6288 1 6286
2 6290 1 6289
2 6291 1 6289
2 6293 1 6292
2 6294 1 6292
2 6296 1 6295
2 6297 1 6295
2 6299 1 6298
2 6300 1 6298
2 6302 1 6301
2 6303 1 6301
2 6305 1 6304
2 6306 1 6304
2 6308 1 6307
2 6309 1 6307
2 6311 1 6310
2 6312 1 6310
2 6314 1 6313
2 6315 1 6313
2 6317 1 6316
2 6318 1 6316
2 6320 1 6319
2 6321 1 6319
2 6323 1 6322
2 6324 1 6322
2 6326 1 6325
2 6327 1 6325
2 6329 1 6328
2 6330 1 6328
2 6332 1 6331
2 6333 1 6331
2 6336 1 6335
2 6337 1 6335
2 6339 1 6338
2 6340 1 6338
2 6342 1 6341
2 6343 1 6341
2 6345 1 6344
2 6346 1 6344
2 6348 1 6347
2 6349 1 6347
2 6351 1 6350
2 6352 1 6350
2 6354 1 6353
2 6355 1 6353
2 6357 1 6356
2 6358 1 6356
2 6360 1 6359
2 6361 1 6359
2 6365 1 6364
2 6366 1 6364
2 6368 1 6367
2 6369 1 6367
2 6371 1 6370
2 6372 1 6370
2 6398 1 6397
2 6399 1 6397
2 6412 1 6411
2 6413 1 6411
2 6416 1 6415
2 6417 1 6415
2 6418 1 6415
2 6420 1 6419
2 6421 1 6419
2 6428 1 6427
2 6429 1 6427
2 6438 1 6437
2 6439 1 6437
2 6442 1 6441
2 6443 1 6441
2 6444 1 6441
2 6446 1 6445
2 6447 1 6445
2 6467 1 6466
2 6468 1 6466
2 6479 1 6478
2 6480 1 6478
2 6483 1 6482
2 6484 1 6482
2 6487 1 6486
2 6488 1 6486
2 6491 1 6490
2 6492 1 6490
2 6495 1 6494
2 6496 1 6494
2 6501 1 6500
2 6502 1 6500
2 6505 1 6504
2 6506 1 6504
2 6509 1 6508
2 6510 1 6508
2 6513 1 6512
2 6514 1 6512
2 6517 1 6516
2 6518 1 6516
2 6527 1 6526
2 6528 1 6526
2 6537 1 6536
2 6538 1 6536
2 6540 1 6539
2 6541 1 6539
2 6554 1 6553
2 6555 1 6553
2 6557 1 6556
2 6558 1 6556
2 6567 1 6566
2 6568 1 6566
2 6570 1 6569
2 6571 1 6569
2 6573 1 6572
2 6574 1 6572
2 6576 1 6575
2 6577 1 6575
2 6581 1 6580
2 6582 1 6580
2 6585 1 6584
2 6586 1 6584
2 6588 1 6587
2 6589 1 6587
2 6593 1 6592
2 6594 1 6592
2 6600 1 6599
2 6601 1 6599
2 6607 1 6606
2 6608 1 6606
2 6610 1 6609
2 6611 1 6609
2 6620 1 6619
2 6621 1 6619
2 6623 1 6622
2 6624 1 6622
2 6635 1 6634
2 6636 1 6634
2 6638 1 6637
2 6639 1 6637
2 6725 1 6724
2 6726 1 6724
2 6793 1 6792
2 6794 1 6792
2 6796 1 6795
2 6797 1 6795
2 6818 1 6817
2 6819 1 6817
2 6820 1 6817
2 6821 1 6817
2 6822 1 6817
2 6832 1 6831
2 6833 1 6831
2 6845 1 6844
2 6846 1 6844
2 6847 1 6844
2 6848 1 6844
2 6849 1 6844
2 6858 1 6857
2 6859 1 6857
2 6867 1 6866
2 6868 1 6866
2 6869 1 6866
2 6870 1 6866
2 6871 1 6866
2 6882 1 6881
2 6883 1 6881
2 6886 1 6885
2 6887 1 6885
2 6892 1 6891
2 6893 1 6891
2 6898 1 6897
2 6899 1 6897
2 6902 1 6901
2 6903 1 6901
2 6906 1 6905
2 6907 1 6905
2 6910 1 6909
2 6911 1 6909
2 6917 1 6916
2 6918 1 6916
2 6933 1 6932
2 6934 1 6932
2 6968 1 6967
2 6969 1 6967
2 6980 1 6979
2 6981 1 6979
2 6982 1 6979
2 7004 1 7003
2 7005 1 7003
2 7007 1 7006
2 7008 1 7006
2 7024 1 7023
2 7025 1 7023
2 7026 1 7023
2 7027 1 7023
2 7029 1 7028
2 7030 1 7028
2 7032 1 7031
2 7033 1 7031
2 7035 1 7034
2 7036 1 7034
2 7038 1 7037
2 7039 1 7037
2 7042 1 7041
2 7043 1 7041
2 7050 1 7049
2 7051 1 7049
2 7052 1 7049
2 7053 1 7049
2 7055 1 7054
2 7056 1 7054
2 7058 1 7057
2 7059 1 7057
2 7061 1 7060
2 7062 1 7060
2 7066 1 7065
2 7067 1 7065
2 7077 1 7076
2 7078 1 7076
2 7081 1 7080
2 7082 1 7080
2 7091 1 7090
2 7092 1 7090
2 7095 1 7094
2 7096 1 7094
2 7098 1 7097
2 7099 1 7097
2 7102 1 7101
2 7103 1 7101
2 7191 1 7190
2 7192 1 7190
2 7193 1 7190
2 7194 1 7190
2 7195 1 7190
2 7199 1 7198
2 7200 1 7198
2 7201 1 7198
2 7202 1 7198
2 7203 1 7198
2 7210 1 7209
2 7211 1 7209
2 7213 1 7212
2 7214 1 7212
2 7220 1 7219
2 7221 1 7219
2 7223 1 7222
2 7224 1 7222
2 7226 1 7225
2 7227 1 7225
2 7237 1 7236
2 7238 1 7236
2 7240 1 7239
2 7241 1 7239
2 7243 1 7242
2 7244 1 7242
2 7246 1 7245
2 7247 1 7245
2 7251 1 7250
2 7252 1 7250
2 7253 1 7250
2 7254 1 7250
2 7255 1 7250
2 7256 1 7250
2 7258 1 7257
2 7259 1 7257
2 7261 1 7260
2 7262 1 7260
2 7264 1 7263
2 7265 1 7263
2 7271 1 7270
2 7272 1 7270
2 7273 1 7270
2 7274 1 7270
2 7275 1 7270
2 7277 1 7276
2 7278 1 7276
2 7279 1 7276
2 7280 1 7276
2 7281 1 7276
2 7283 1 7282
2 7284 1 7282
2 7285 1 7282
2 7286 1 7282
2 7287 1 7282
2 7289 1 7288
2 7290 1 7288
2 7291 1 7288
2 7292 1 7288
2 7293 1 7288
2 7295 1 7294
2 7296 1 7294
2 7297 1 7294
2 7298 1 7294
2 7299 1 7294
2 7302 1 7301
2 7303 1 7301
2 7305 1 7304
2 7306 1 7304
2 7307 1 7304
2 7308 1 7304
2 7309 1 7304
2 7311 1 7310
2 7312 1 7310
2 7313 1 7310
2 7314 1 7310
2 7315 1 7310
2 7395 1 7394
2 7396 1 7394
2 7398 1 7397
2 7399 1 7397
2 7403 1 7402
2 7404 1 7402
2 7410 1 7409
2 7411 1 7409
2 7413 1 7412
2 7414 1 7412
2 7422 1 7421
2 7423 1 7421
2 7490 1 7489
2 7491 1 7489
2 7532 1 7531
2 7533 1 7531
2 7534 1 7531
2 7535 1 7531
2 7536 1 7531
2 7538 1 7537
2 7539 1 7537
2 7540 1 7537
2 7541 1 7537
2 7542 1 7537
2 7544 1 7543
2 7545 1 7543
2 7546 1 7543
2 7547 1 7543
2 7548 1 7543
2 7550 1 7549
2 7551 1 7549
2 7552 1 7549
2 7553 1 7549
2 7554 1 7549
2 7556 1 7555
2 7557 1 7555
2 7558 1 7555
2 7559 1 7555
2 7560 1 7555
2 7562 1 7561
2 7563 1 7561
2 7564 1 7561
2 7565 1 7561
2 7566 1 7561
2 7568 1 7567
2 7569 1 7567
2 7570 1 7567
2 7571 1 7567
2 7572 1 7567
2 7574 1 7573
2 7575 1 7573
2 7576 1 7573
2 7577 1 7573
2 7578 1 7573
2 7580 1 7579
2 7581 1 7579
2 7583 1 7582
2 7584 1 7582
2 7590 1 7589
2 7591 1 7589
2 7593 1 7592
2 7594 1 7592
2 7596 1 7595
2 7597 1 7595
2 7713 1 7712
2 7714 1 7712
2 7716 1 7715
2 7717 1 7715
2 7725 1 7724
2 7726 1 7724
2 7763 1 7762
2 7764 1 7762
2 7766 1 7765
2 7767 1 7765
2 7773 1 7772
2 7774 1 7772
2 7776 1 7775
2 7777 1 7775
2 7779 1 7778
2 7780 1 7778
2 7801 1 7800
2 7802 1 7800
2 7804 1 7803
2 7805 1 7803
2 7813 1 7812
2 7814 1 7812
2 7827 1 7826
2 7828 1 7826
2 7830 1 7829
2 7831 1 7829
2 7837 1 7836
2 7838 1 7836
2 7840 1 7839
2 7841 1 7839
2 7843 1 7842
2 7844 1 7842
2 7865 1 7864
2 7866 1 7864
2 7868 1 7867
2 7869 1 7867
2 7877 1 7876
2 7878 1 7876
2 7891 1 7890
2 7892 1 7890
2 7894 1 7893
2 7895 1 7893
2 7901 1 7900
2 7902 1 7900
2 7904 1 7903
2 7905 1 7903
2 7907 1 7906
2 7908 1 7906
2 7933 1 7932
2 7934 1 7932
2 7936 1 7935
2 7937 1 7935
2 7941 1 7940
2 7942 1 7940
2 7955 1 7954
2 7956 1 7954
2 7958 1 7957
2 7959 1 7957
2 7961 1 7960
2 7962 1 7960
2 7964 1 7963
2 7965 1 7963
2 7971 1 7970
2 7972 1 7970
2 7999 1 7998
2 8000 1 7998
2 8002 1 8001
2 8003 1 8001
2 8005 1 8004
2 8006 1 8004
2 8014 1 8013
2 8015 1 8013
2 8018 1 8017
2 8019 1 8017
2 8046 1 8045
2 8047 1 8045
2 8049 1 8048
2 8050 1 8048
2 8062 1 8061
2 8063 1 8061
2 8065 1 8064
2 8066 1 8064
2 8080 1 8079
2 8081 1 8079
2 8083 1 8082
2 8084 1 8082
2 8094 1 8093
2 8095 1 8093
2 8097 1 8096
2 8098 1 8096
2 8100 1 8099
2 8101 1 8099
2 8103 1 8102
2 8104 1 8102
